/*
 * This file is automatically generated
 * k = 4, M = 8
 */ 

module crossbar (
  input clk,    // Clock
  input clk_en, // Clock Enable
  input in0,input in1,input in2,
);

  assign out0 = in0;

  always@(posedge clk) begin
    if (clk_en) begin
      out0_reg <= out0;


endmodule