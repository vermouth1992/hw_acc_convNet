// Latency: 31
// Gap: 1
module codeBlock22226(clk, reset, next_in, next_out,
   X0_in, Y0,
   X1_in, Y1,
   X2_in, Y2,
   X3_in, Y3,
   X4_in, Y4,
   X5_in, Y5,
   X6_in, Y6,
   X7_in, Y7,
   X8_in, Y8,
   X9_in, Y9,
   X10_in, Y10,
   X11_in, Y11,
   X12_in, Y12,
   X13_in, Y13,
   X14_in, Y14,
   X15_in, Y15);

   output next_out;
   input clk, reset, next_in;

   reg next;

   input [31:0] X0_in,
      X1_in,
      X2_in,
      X3_in,
      X4_in,
      X5_in,
      X6_in,
      X7_in,
      X8_in,
      X9_in,
      X10_in,
      X11_in,
      X12_in,
      X13_in,
      X14_in,
      X15_in;

   reg   [31:0] X0,
      X1,
      X2,
      X3,
      X4,
      X5,
      X6,
      X7,
      X8,
      X9,
      X10,
      X11,
      X12,
      X13,
      X14,
      X15;

   output [31:0] Y0,
      Y1,
      Y2,
      Y3,
      Y4,
      Y5,
      Y6,
      Y7,
      Y8,
      Y9,
      Y10,
      Y11,
      Y12,
      Y13,
      Y14,
      Y15;

   shiftRegFIFO #(30, 1) shiftFIFO_23923(.X(next), .Y(next_out), .clk(clk));


   wire signed [31:0] a109;
   wire signed [31:0] a110;
   wire signed [31:0] a111;
   wire signed [31:0] a112;
   wire signed [31:0] a117;
   wire signed [31:0] a118;
   wire signed [31:0] a119;
   wire signed [31:0] a120;
   wire signed [31:0] a125;
   wire signed [31:0] a126;
   wire signed [31:0] a127;
   wire signed [31:0] a128;
   wire signed [31:0] a133;
   wire signed [31:0] a134;
   wire signed [31:0] a135;
   wire signed [31:0] a136;
   wire  [31:0] t349;
   wire  [31:0] t350;
   wire  [31:0] t351;
   wire  [31:0] t352;
   wire  [31:0] t353;
   wire  [31:0] t354;
   wire  [31:0] t355;
   wire  [31:0] t356;
   wire  [31:0] t359;
   wire  [31:0] t360;
   wire  [31:0] t361;
   wire  [31:0] t362;
   wire  [31:0] t363;
   wire  [31:0] t364;
   wire  [31:0] t365;
   wire  [31:0] t366;
   reg signed [31:0] tm4;
   reg signed [31:0] tm23;
   reg signed [31:0] tm42;
   reg signed [31:0] tm61;
   reg signed [31:0] tm80;
   reg signed [31:0] tm99;
   reg signed [31:0] tm118;
   reg signed [31:0] tm137;
   reg signed [31:0] tm156;
   reg signed [31:0] tm175;
   reg signed [31:0] tm194;
   reg signed [31:0] tm213;
   reg signed [31:0] tm5;
   reg signed [31:0] tm24;
   reg signed [31:0] tm43;
   reg signed [31:0] tm62;
   reg signed [31:0] tm81;
   reg signed [31:0] tm100;
   reg signed [31:0] tm119;
   reg signed [31:0] tm138;
   reg signed [31:0] tm157;
   reg signed [31:0] tm176;
   reg signed [31:0] tm195;
   reg signed [31:0] tm214;
   reg signed [31:0] tm6;
   reg signed [31:0] tm25;
   reg signed [31:0] tm44;
   reg signed [31:0] tm63;
   reg signed [31:0] tm82;
   reg signed [31:0] tm101;
   reg signed [31:0] tm120;
   reg signed [31:0] tm139;
   reg signed [31:0] tm158;
   reg signed [31:0] tm177;
   reg signed [31:0] tm196;
   reg signed [31:0] tm215;
   reg signed [31:0] tm7;
   reg signed [31:0] tm26;
   reg signed [31:0] tm45;
   reg signed [31:0] tm64;
   reg signed [31:0] tm83;
   reg signed [31:0] tm102;
   reg signed [31:0] tm121;
   reg signed [31:0] tm140;
   reg signed [31:0] tm159;
   reg signed [31:0] tm178;
   reg signed [31:0] tm197;
   reg signed [31:0] tm216;
   reg signed [31:0] tm8;
   reg signed [31:0] tm27;
   reg signed [31:0] tm46;
   reg signed [31:0] tm65;
   reg signed [31:0] tm84;
   reg signed [31:0] tm103;
   reg signed [31:0] tm122;
   reg signed [31:0] tm141;
   reg signed [31:0] tm160;
   reg signed [31:0] tm179;
   reg signed [31:0] tm198;
   reg signed [31:0] tm217;
   reg signed [31:0] tm9;
   reg signed [31:0] tm28;
   reg signed [31:0] tm47;
   reg signed [31:0] tm66;
   reg signed [31:0] tm85;
   reg signed [31:0] tm104;
   reg signed [31:0] tm123;
   reg signed [31:0] tm142;
   reg signed [31:0] tm161;
   reg signed [31:0] tm180;
   reg signed [31:0] tm199;
   reg signed [31:0] tm218;
   reg signed [31:0] tm10;
   reg signed [31:0] tm29;
   reg signed [31:0] tm48;
   reg signed [31:0] tm67;
   reg signed [31:0] tm86;
   reg signed [31:0] tm105;
   reg signed [31:0] tm124;
   reg signed [31:0] tm143;
   reg signed [31:0] tm162;
   reg signed [31:0] tm181;
   reg signed [31:0] tm200;
   reg signed [31:0] tm219;
   wire  [31:0] a105;
   wire  [31:0] a106;
   wire  [31:0] a107;
   wire  [31:0] a108;
   reg signed [31:0] tm11;
   reg signed [31:0] tm30;
   reg signed [31:0] tm49;
   reg signed [31:0] tm68;
   reg signed [31:0] tm87;
   reg signed [31:0] tm106;
   reg signed [31:0] tm125;
   reg signed [31:0] tm144;
   reg signed [31:0] tm163;
   reg signed [31:0] tm182;
   reg signed [31:0] tm201;
   reg signed [31:0] tm220;
   reg signed [31:0] tm12;
   reg signed [31:0] tm31;
   reg signed [31:0] tm50;
   reg signed [31:0] tm69;
   reg signed [31:0] tm88;
   reg signed [31:0] tm107;
   reg signed [31:0] tm126;
   reg signed [31:0] tm145;
   reg signed [31:0] tm164;
   reg signed [31:0] tm183;
   reg signed [31:0] tm202;
   reg signed [31:0] tm221;
   reg signed [31:0] tm13;
   reg signed [31:0] tm32;
   reg signed [31:0] tm51;
   reg signed [31:0] tm70;
   reg signed [31:0] tm89;
   reg signed [31:0] tm108;
   reg signed [31:0] tm127;
   reg signed [31:0] tm146;
   reg signed [31:0] tm165;
   reg signed [31:0] tm184;
   reg signed [31:0] tm203;
   reg signed [31:0] tm222;
   reg signed [31:0] tm14;
   reg signed [31:0] tm33;
   reg signed [31:0] tm52;
   reg signed [31:0] tm71;
   reg signed [31:0] tm90;
   reg signed [31:0] tm109;
   reg signed [31:0] tm128;
   reg signed [31:0] tm147;
   reg signed [31:0] tm166;
   reg signed [31:0] tm185;
   reg signed [31:0] tm204;
   reg signed [31:0] tm223;
   reg signed [31:0] tm15;
   reg signed [31:0] tm34;
   reg signed [31:0] tm53;
   reg signed [31:0] tm72;
   reg signed [31:0] tm91;
   reg signed [31:0] tm110;
   reg signed [31:0] tm129;
   reg signed [31:0] tm148;
   reg signed [31:0] tm167;
   reg signed [31:0] tm186;
   reg signed [31:0] tm205;
   reg signed [31:0] tm224;
   reg signed [31:0] tm16;
   reg signed [31:0] tm35;
   reg signed [31:0] tm54;
   reg signed [31:0] tm73;
   reg signed [31:0] tm92;
   reg signed [31:0] tm111;
   reg signed [31:0] tm130;
   reg signed [31:0] tm149;
   reg signed [31:0] tm168;
   reg signed [31:0] tm187;
   reg signed [31:0] tm206;
   reg signed [31:0] tm225;
   reg signed [31:0] tm17;
   reg signed [31:0] tm36;
   reg signed [31:0] tm55;
   reg signed [31:0] tm74;
   reg signed [31:0] tm93;
   reg signed [31:0] tm112;
   reg signed [31:0] tm131;
   reg signed [31:0] tm150;
   reg signed [31:0] tm169;
   reg signed [31:0] tm188;
   reg signed [31:0] tm207;
   reg signed [31:0] tm226;
   reg signed [31:0] tm18;
   reg signed [31:0] tm37;
   reg signed [31:0] tm56;
   reg signed [31:0] tm75;
   reg signed [31:0] tm94;
   reg signed [31:0] tm113;
   reg signed [31:0] tm132;
   reg signed [31:0] tm151;
   reg signed [31:0] tm170;
   reg signed [31:0] tm189;
   reg signed [31:0] tm208;
   reg signed [31:0] tm227;
   reg signed [31:0] tm19;
   reg signed [31:0] tm38;
   reg signed [31:0] tm57;
   reg signed [31:0] tm76;
   reg signed [31:0] tm95;
   reg signed [31:0] tm114;
   reg signed [31:0] tm133;
   reg signed [31:0] tm152;
   reg signed [31:0] tm171;
   reg signed [31:0] tm190;
   reg signed [31:0] tm209;
   reg signed [31:0] tm228;
   reg signed [31:0] tm20;
   reg signed [31:0] tm39;
   reg signed [31:0] tm58;
   reg signed [31:0] tm77;
   reg signed [31:0] tm96;
   reg signed [31:0] tm115;
   reg signed [31:0] tm134;
   reg signed [31:0] tm153;
   reg signed [31:0] tm172;
   reg signed [31:0] tm191;
   reg signed [31:0] tm210;
   reg signed [31:0] tm229;
   reg signed [31:0] tm21;
   reg signed [31:0] tm40;
   reg signed [31:0] tm59;
   reg signed [31:0] tm78;
   reg signed [31:0] tm97;
   reg signed [31:0] tm116;
   reg signed [31:0] tm135;
   reg signed [31:0] tm154;
   reg signed [31:0] tm173;
   reg signed [31:0] tm192;
   reg signed [31:0] tm211;
   reg signed [31:0] tm230;
   wire signed [31:0] Y0;
   wire signed [31:0] Y1;
   wire signed [31:0] Y2;
   wire signed [31:0] Y3;
   wire  [31:0] t357;
   wire  [31:0] t358;
   wire signed [31:0] Y4;
   wire signed [31:0] Y5;
   wire signed [31:0] Y6;
   wire signed [31:0] Y7;
   wire signed [31:0] Y8;
   wire signed [31:0] Y9;
   wire signed [31:0] Y10;
   wire signed [31:0] Y11;
   wire  [31:0] t367;
   wire  [31:0] t368;
   wire signed [31:0] Y12;
   wire signed [31:0] Y13;
   wire signed [31:0] Y14;
   wire signed [31:0] Y15;
   reg signed [31:0] tm22;
   reg signed [31:0] tm41;
   reg signed [31:0] tm60;
   reg signed [31:0] tm79;
   reg signed [31:0] tm98;
   reg signed [31:0] tm117;
   reg signed [31:0] tm136;
   reg signed [31:0] tm155;
   reg signed [31:0] tm174;
   reg signed [31:0] tm193;
   reg signed [31:0] tm212;
   reg signed [31:0] tm231;

   wire signed [31:0] tm0;
   assign tm0 = 32'h3f3504f3;

   assign a109 = X0;
   assign a110 = X8;
   assign a111 = X1;
   assign a112 = X9;
   assign a117 = X2;
   assign a118 = X10;
   assign a119 = X3;
   assign a120 = X11;
   assign a125 = X4;
   assign a126 = X12;
   assign a127 = X5;
   assign a128 = X13;
   assign a133 = X6;
   assign a134 = X14;
   assign a135 = X7;
   assign a136 = X15;
   assign Y0 = tm22;
   assign Y1 = tm41;
   assign Y2 = tm60;
   assign Y3 = tm79;
   assign Y4 = tm98;
   assign Y5 = tm117;
   assign Y6 = t357;
   assign Y7 = t358;
   assign Y8 = tm136;
   assign Y9 = tm155;
   assign Y10 = tm174;
   assign Y11 = tm193;
   assign Y12 = tm212;
   assign Y13 = tm231;
   assign Y14 = {~(t367[31]), t367[30:0]};
   assign Y15 = t368;

    addfp32 add22238(.a(a109), .b(a110), .clk(clk), .out(t349), .enable(1'b1), .rst(reset));
    addfp32 add22253(.a(a111), .b(a112), .clk(clk), .out(t350), .enable(1'b1), .rst(reset));
    subfp32 sub22268(.a(a109), .b(a110), .clk(clk), .out(t351), .enable(1'b1), .rst(reset));
    subfp32 sub22283(.a(a111), .b(a112), .clk(clk), .out(t352), .enable(1'b1), .rst(reset));
    addfp32 add22314(.a(a117), .b(a118), .clk(clk), .out(t353), .enable(1'b1), .rst(reset));
    addfp32 add22329(.a(a119), .b(a120), .clk(clk), .out(t354), .enable(1'b1), .rst(reset));
    subfp32 sub22344(.a(a117), .b(a118), .clk(clk), .out(t355), .enable(1'b1), .rst(reset));
    subfp32 sub22359(.a(a119), .b(a120), .clk(clk), .out(t356), .enable(1'b1), .rst(reset));
    addfp32 add22418(.a(a125), .b(a126), .clk(clk), .out(t359), .enable(1'b1), .rst(reset));
    addfp32 add22433(.a(a127), .b(a128), .clk(clk), .out(t360), .enable(1'b1), .rst(reset));
    subfp32 sub22448(.a(a125), .b(a126), .clk(clk), .out(t361), .enable(1'b1), .rst(reset));
    subfp32 sub22463(.a(a127), .b(a128), .clk(clk), .out(t362), .enable(1'b1), .rst(reset));
    addfp32 add22495(.a(a133), .b(a134), .clk(clk), .out(t363), .enable(1'b1), .rst(reset));
    addfp32 add22510(.a(a135), .b(a136), .clk(clk), .out(t364), .enable(1'b1), .rst(reset));
    subfp32 sub22525(.a(a133), .b(a134), .clk(clk), .out(t365), .enable(1'b1), .rst(reset));
    subfp32 sub22540(.a(a135), .b(a136), .clk(clk), .out(t366), .enable(1'b1), .rst(reset));
    multfp32fp32 m22366(.a(tm0), .b(t355), .clk(clk), .out(a105), .enable(1'b1), .rst(reset));
    multfp32fp32 m22373(.a(tm0), .b(t356), .clk(clk), .out(a106), .enable(1'b1), .rst(reset));
    multfp32fp32 m22547(.a(tm0), .b(t365), .clk(clk), .out(a107), .enable(1'b1), .rst(reset));
    multfp32fp32 m22554(.a(tm0), .b(t366), .clk(clk), .out(a108), .enable(1'b1), .rst(reset));
    subfp32 sub22380(.a(a105), .b(a106), .clk(clk), .out(t357), .enable(1'b1), .rst(reset));
    addfp32 add22387(.a(a105), .b(a106), .clk(clk), .out(t358), .enable(1'b1), .rst(reset));
    addfp32 add22561(.a(a107), .b(a108), .clk(clk), .out(t367), .enable(1'b1), .rst(reset));
    subfp32 sub22568(.a(a107), .b(a108), .clk(clk), .out(t368), .enable(1'b1), .rst(reset));


   always @(posedge clk) begin
      if (reset == 1) begin
      end
      else begin
         X0 <= X0_in;
         X1 <= X1_in;
         X2 <= X2_in;
         X3 <= X3_in;
         X4 <= X4_in;
         X5 <= X5_in;
         X6 <= X6_in;
         X7 <= X7_in;
         X8 <= X8_in;
         X9 <= X9_in;
         X10 <= X10_in;
         X11 <= X11_in;
         X12 <= X12_in;
         X13 <= X13_in;
         X14 <= X14_in;
         X15 <= X15_in;
         next <= next_in;
         tm4 <= t349;
         tm23 <= t350;
         tm42 <= t351;
         tm61 <= t352;
         tm80 <= t353;
         tm99 <= t354;
         tm118 <= t359;
         tm137 <= t360;
         tm156 <= {~(t362[31]), t362[30:0]};
         tm175 <= t361;
         tm194 <= t363;
         tm213 <= t364;
         tm5 <= tm4;
         tm24 <= tm23;
         tm43 <= tm42;
         tm62 <= tm61;
         tm81 <= tm80;
         tm100 <= tm99;
         tm119 <= tm118;
         tm138 <= tm137;
         tm157 <= tm156;
         tm176 <= tm175;
         tm195 <= tm194;
         tm214 <= tm213;
         tm6 <= tm5;
         tm25 <= tm24;
         tm44 <= tm43;
         tm63 <= tm62;
         tm82 <= tm81;
         tm101 <= tm100;
         tm120 <= tm119;
         tm139 <= tm138;
         tm158 <= tm157;
         tm177 <= tm176;
         tm196 <= tm195;
         tm215 <= tm214;
         tm7 <= tm6;
         tm26 <= tm25;
         tm45 <= tm44;
         tm64 <= tm63;
         tm83 <= tm82;
         tm102 <= tm101;
         tm121 <= tm120;
         tm140 <= tm139;
         tm159 <= tm158;
         tm178 <= tm177;
         tm197 <= tm196;
         tm216 <= tm215;
         tm8 <= tm7;
         tm27 <= tm26;
         tm46 <= tm45;
         tm65 <= tm64;
         tm84 <= tm83;
         tm103 <= tm102;
         tm122 <= tm121;
         tm141 <= tm140;
         tm160 <= tm159;
         tm179 <= tm178;
         tm198 <= tm197;
         tm217 <= tm216;
         tm9 <= tm8;
         tm28 <= tm27;
         tm47 <= tm46;
         tm66 <= tm65;
         tm85 <= tm84;
         tm104 <= tm103;
         tm123 <= tm122;
         tm142 <= tm141;
         tm161 <= tm160;
         tm180 <= tm179;
         tm199 <= tm198;
         tm218 <= tm217;
         tm10 <= tm9;
         tm29 <= tm28;
         tm48 <= tm47;
         tm67 <= tm66;
         tm86 <= tm85;
         tm105 <= tm104;
         tm124 <= tm123;
         tm143 <= tm142;
         tm162 <= tm161;
         tm181 <= tm180;
         tm200 <= tm199;
         tm219 <= tm218;
         tm11 <= tm10;
         tm30 <= tm29;
         tm49 <= tm48;
         tm68 <= tm67;
         tm87 <= tm86;
         tm106 <= tm105;
         tm125 <= tm124;
         tm144 <= tm143;
         tm163 <= tm162;
         tm182 <= tm181;
         tm201 <= tm200;
         tm220 <= tm219;
         tm12 <= tm11;
         tm31 <= tm30;
         tm50 <= tm49;
         tm69 <= tm68;
         tm88 <= tm87;
         tm107 <= tm106;
         tm126 <= tm125;
         tm145 <= tm144;
         tm164 <= tm163;
         tm183 <= tm182;
         tm202 <= tm201;
         tm221 <= tm220;
         tm13 <= tm12;
         tm32 <= tm31;
         tm51 <= tm50;
         tm70 <= tm69;
         tm89 <= tm88;
         tm108 <= tm107;
         tm127 <= tm126;
         tm146 <= tm145;
         tm165 <= tm164;
         tm184 <= tm183;
         tm203 <= tm202;
         tm222 <= tm221;
         tm14 <= tm13;
         tm33 <= tm32;
         tm52 <= tm51;
         tm71 <= tm70;
         tm90 <= tm89;
         tm109 <= tm108;
         tm128 <= tm127;
         tm147 <= tm146;
         tm166 <= tm165;
         tm185 <= tm184;
         tm204 <= tm203;
         tm223 <= tm222;
         tm15 <= tm14;
         tm34 <= tm33;
         tm53 <= tm52;
         tm72 <= tm71;
         tm91 <= tm90;
         tm110 <= tm109;
         tm129 <= tm128;
         tm148 <= tm147;
         tm167 <= tm166;
         tm186 <= tm185;
         tm205 <= tm204;
         tm224 <= tm223;
         tm16 <= tm15;
         tm35 <= tm34;
         tm54 <= tm53;
         tm73 <= tm72;
         tm92 <= tm91;
         tm111 <= tm110;
         tm130 <= tm129;
         tm149 <= tm148;
         tm168 <= tm167;
         tm187 <= tm186;
         tm206 <= tm205;
         tm225 <= tm224;
         tm17 <= tm16;
         tm36 <= tm35;
         tm55 <= tm54;
         tm74 <= tm73;
         tm93 <= tm92;
         tm112 <= tm111;
         tm131 <= tm130;
         tm150 <= tm149;
         tm169 <= tm168;
         tm188 <= tm187;
         tm207 <= tm206;
         tm226 <= tm225;
         tm18 <= tm17;
         tm37 <= tm36;
         tm56 <= tm55;
         tm75 <= tm74;
         tm94 <= tm93;
         tm113 <= tm112;
         tm132 <= tm131;
         tm151 <= tm150;
         tm170 <= tm169;
         tm189 <= tm188;
         tm208 <= tm207;
         tm227 <= tm226;
         tm19 <= tm18;
         tm38 <= tm37;
         tm57 <= tm56;
         tm76 <= tm75;
         tm95 <= tm94;
         tm114 <= tm113;
         tm133 <= tm132;
         tm152 <= tm151;
         tm171 <= tm170;
         tm190 <= tm189;
         tm209 <= tm208;
         tm228 <= tm227;
         tm20 <= tm19;
         tm39 <= tm38;
         tm58 <= tm57;
         tm77 <= tm76;
         tm96 <= tm95;
         tm115 <= tm114;
         tm134 <= tm133;
         tm153 <= tm152;
         tm172 <= tm171;
         tm191 <= tm190;
         tm210 <= tm209;
         tm229 <= tm228;
         tm21 <= tm20;
         tm40 <= tm39;
         tm59 <= tm58;
         tm78 <= tm77;
         tm97 <= tm96;
         tm116 <= tm115;
         tm135 <= tm134;
         tm154 <= tm153;
         tm173 <= tm172;
         tm192 <= tm191;
         tm211 <= tm210;
         tm230 <= tm229;
         tm22 <= tm21;
         tm41 <= tm40;
         tm60 <= tm59;
         tm79 <= tm78;
         tm98 <= tm97;
         tm117 <= tm116;
         tm136 <= tm135;
         tm155 <= tm154;
         tm174 <= tm173;
         tm193 <= tm192;
         tm212 <= tm211;
         tm231 <= tm230;
      end
   end
endmodule

// Latency: 23
// Gap: 1
module codeBlock22590(clk, reset, next_in, next_out,
   X0_in, Y0,
   X1_in, Y1,
   X2_in, Y2,
   X3_in, Y3,
   X4_in, Y4,
   X5_in, Y5,
   X6_in, Y6,
   X7_in, Y7,
   X8_in, Y8,
   X9_in, Y9,
   X10_in, Y10,
   X11_in, Y11,
   X12_in, Y12,
   X13_in, Y13,
   X14_in, Y14,
   X15_in, Y15);

   output next_out;
   input clk, reset, next_in;

   reg next;

   input [31:0] X0_in,
      X1_in,
      X2_in,
      X3_in,
      X4_in,
      X5_in,
      X6_in,
      X7_in,
      X8_in,
      X9_in,
      X10_in,
      X11_in,
      X12_in,
      X13_in,
      X14_in,
      X15_in;

   reg   [31:0] X0,
      X1,
      X2,
      X3,
      X4,
      X5,
      X6,
      X7,
      X8,
      X9,
      X10,
      X11,
      X12,
      X13,
      X14,
      X15;

   output [31:0] Y0,
      Y1,
      Y2,
      Y3,
      Y4,
      Y5,
      Y6,
      Y7,
      Y8,
      Y9,
      Y10,
      Y11,
      Y12,
      Y13,
      Y14,
      Y15;

   shiftRegFIFO #(22, 1) shiftFIFO_23926(.X(next), .Y(next_out), .clk(clk));


   wire signed [31:0] a33;
   wire signed [31:0] a34;
   wire signed [31:0] a35;
   wire signed [31:0] a36;
   wire signed [31:0] a41;
   wire signed [31:0] a42;
   wire signed [31:0] a43;
   wire signed [31:0] a44;
   wire signed [31:0] a49;
   wire signed [31:0] a50;
   wire signed [31:0] a51;
   wire signed [31:0] a52;
   wire signed [31:0] a57;
   wire signed [31:0] a58;
   wire signed [31:0] a59;
   wire signed [31:0] a60;
   wire  [31:0] t209;
   wire  [31:0] t210;
   wire  [31:0] t211;
   wire  [31:0] t212;
   wire  [31:0] t213;
   wire  [31:0] t214;
   wire  [31:0] t215;
   wire  [31:0] t216;
   wire  [31:0] t225;
   wire  [31:0] t226;
   wire  [31:0] t227;
   wire  [31:0] t228;
   wire  [31:0] t229;
   wire  [31:0] t230;
   wire  [31:0] t231;
   wire  [31:0] t232;
   wire  [31:0] t217;
   wire  [31:0] t218;
   wire  [31:0] t219;
   wire  [31:0] t220;
   wire signed [31:0] Y0;
   wire signed [31:0] Y1;
   wire signed [31:0] Y8;
   wire signed [31:0] Y9;
   wire  [31:0] t221;
   wire  [31:0] t222;
   wire  [31:0] t223;
   wire  [31:0] t224;
   wire signed [31:0] Y4;
   wire signed [31:0] Y5;
   wire signed [31:0] Y12;
   wire signed [31:0] Y13;
   wire  [31:0] t233;
   wire  [31:0] t234;
   wire  [31:0] t235;
   wire  [31:0] t236;
   wire signed [31:0] Y2;
   wire signed [31:0] Y3;
   wire signed [31:0] Y10;
   wire signed [31:0] Y11;
   wire  [31:0] t237;
   wire  [31:0] t238;
   wire  [31:0] t239;
   wire  [31:0] t240;
   wire signed [31:0] Y6;
   wire signed [31:0] Y7;
   wire signed [31:0] Y14;
   wire signed [31:0] Y15;


   assign a33 = X0;
   assign a34 = X8;
   assign a35 = X1;
   assign a36 = X9;
   assign a41 = X4;
   assign a42 = X12;
   assign a43 = X5;
   assign a44 = X13;
   assign a49 = X2;
   assign a50 = X10;
   assign a51 = X3;
   assign a52 = X11;
   assign a57 = X6;
   assign a58 = X14;
   assign a59 = X7;
   assign a60 = X15;
   assign Y0 = t217;
   assign Y1 = t218;
   assign Y8 = t219;
   assign Y9 = t220;
   assign Y4 = t221;
   assign Y5 = t222;
   assign Y12 = t223;
   assign Y13 = t224;
   assign Y2 = t233;
   assign Y3 = t234;
   assign Y10 = t235;
   assign Y11 = t236;
   assign Y6 = t237;
   assign Y7 = t238;
   assign Y14 = t239;
   assign Y15 = t240;

    addfp32 add22602(.a(a33), .b(a34), .clk(clk), .out(t209), .enable(1'b1), .rst(reset));
    addfp32 add22617(.a(a35), .b(a36), .clk(clk), .out(t210), .enable(1'b1), .rst(reset));
    subfp32 sub22632(.a(a33), .b(a34), .clk(clk), .out(t211), .enable(1'b1), .rst(reset));
    subfp32 sub22647(.a(a35), .b(a36), .clk(clk), .out(t212), .enable(1'b1), .rst(reset));
    addfp32 add22662(.a(a41), .b(a42), .clk(clk), .out(t213), .enable(1'b1), .rst(reset));
    addfp32 add22677(.a(a43), .b(a44), .clk(clk), .out(t214), .enable(1'b1), .rst(reset));
    subfp32 sub22692(.a(a41), .b(a42), .clk(clk), .out(t215), .enable(1'b1), .rst(reset));
    subfp32 sub22707(.a(a43), .b(a44), .clk(clk), .out(t216), .enable(1'b1), .rst(reset));
    addfp32 add22810(.a(a49), .b(a50), .clk(clk), .out(t225), .enable(1'b1), .rst(reset));
    addfp32 add22825(.a(a51), .b(a52), .clk(clk), .out(t226), .enable(1'b1), .rst(reset));
    subfp32 sub22840(.a(a49), .b(a50), .clk(clk), .out(t227), .enable(1'b1), .rst(reset));
    subfp32 sub22855(.a(a51), .b(a52), .clk(clk), .out(t228), .enable(1'b1), .rst(reset));
    addfp32 add22870(.a(a57), .b(a58), .clk(clk), .out(t229), .enable(1'b1), .rst(reset));
    addfp32 add22885(.a(a59), .b(a60), .clk(clk), .out(t230), .enable(1'b1), .rst(reset));
    subfp32 sub22900(.a(a57), .b(a58), .clk(clk), .out(t231), .enable(1'b1), .rst(reset));
    subfp32 sub22915(.a(a59), .b(a60), .clk(clk), .out(t232), .enable(1'b1), .rst(reset));
    addfp32 add22714(.a(t209), .b(t213), .clk(clk), .out(t217), .enable(1'b1), .rst(reset));
    addfp32 add22721(.a(t210), .b(t214), .clk(clk), .out(t218), .enable(1'b1), .rst(reset));
    subfp32 sub22728(.a(t209), .b(t213), .clk(clk), .out(t219), .enable(1'b1), .rst(reset));
    subfp32 sub22735(.a(t210), .b(t214), .clk(clk), .out(t220), .enable(1'b1), .rst(reset));
    subfp32 sub22758(.a(t211), .b(t216), .clk(clk), .out(t221), .enable(1'b1), .rst(reset));
    addfp32 add22765(.a(t212), .b(t215), .clk(clk), .out(t222), .enable(1'b1), .rst(reset));
    addfp32 add22772(.a(t211), .b(t216), .clk(clk), .out(t223), .enable(1'b1), .rst(reset));
    subfp32 sub22779(.a(t212), .b(t215), .clk(clk), .out(t224), .enable(1'b1), .rst(reset));
    addfp32 add22922(.a(t225), .b(t229), .clk(clk), .out(t233), .enable(1'b1), .rst(reset));
    addfp32 add22929(.a(t226), .b(t230), .clk(clk), .out(t234), .enable(1'b1), .rst(reset));
    subfp32 sub22936(.a(t225), .b(t229), .clk(clk), .out(t235), .enable(1'b1), .rst(reset));
    subfp32 sub22943(.a(t226), .b(t230), .clk(clk), .out(t236), .enable(1'b1), .rst(reset));
    subfp32 sub22966(.a(t227), .b(t232), .clk(clk), .out(t237), .enable(1'b1), .rst(reset));
    addfp32 add22973(.a(t228), .b(t231), .clk(clk), .out(t238), .enable(1'b1), .rst(reset));
    addfp32 add22980(.a(t227), .b(t232), .clk(clk), .out(t239), .enable(1'b1), .rst(reset));
    subfp32 sub22987(.a(t228), .b(t231), .clk(clk), .out(t240), .enable(1'b1), .rst(reset));


   always @(posedge clk) begin
      if (reset == 1) begin
      end
      else begin
         X0 <= X0_in;
         X1 <= X1_in;
         X2 <= X2_in;
         X3 <= X3_in;
         X4 <= X4_in;
         X5 <= X5_in;
         X6 <= X6_in;
         X7 <= X7_in;
         X8 <= X8_in;
         X9 <= X9_in;
         X10 <= X10_in;
         X11 <= X11_in;
         X12 <= X12_in;
         X13 <= X13_in;
         X14 <= X14_in;
         X15 <= X15_in;
         next <= next_in;
      end
   end
endmodule

