module crossbar(input clk, input reset,
    input  io_clk_en,
    input  io_start,
    output io_start_next_stage,
    input [63:0] io_in_15,
    input [63:0] io_in_14,
    input [63:0] io_in_13,
    input [63:0] io_in_12,
    input [63:0] io_in_11,
    input [63:0] io_in_10,
    input [63:0] io_in_9,
    input [63:0] io_in_8,
    input [63:0] io_in_7,
    input [63:0] io_in_6,
    input [63:0] io_in_5,
    input [63:0] io_in_4,
    input [63:0] io_in_3,
    input [63:0] io_in_2,
    input [63:0] io_in_1,
    input [63:0] io_in_0,
    output[63:0] io_out_15,
    output[63:0] io_out_14,
    output[63:0] io_out_13,
    output[63:0] io_out_12,
    output[63:0] io_out_11,
    output[63:0] io_out_10,
    output[63:0] io_out_9,
    output[63:0] io_out_8,
    output[63:0] io_out_7,
    output[63:0] io_out_6,
    output[63:0] io_out_5,
    output[63:0] io_out_4,
    output[63:0] io_out_3,
    output[63:0] io_out_2,
    output[63:0] io_out_1,
    output[63:0] io_out_0
);

  reg [63:0] out_reg_0;
  wire[63:0] T0;
  wire T1;
  reg [63:0] out_reg_1;
  wire[63:0] T2;
  reg [63:0] out_reg_2;
  wire[63:0] T3;
  reg [63:0] out_reg_3;
  wire[63:0] T4;
  reg [63:0] out_reg_4;
  wire[63:0] T5;
  reg [63:0] out_reg_5;
  wire[63:0] T6;
  reg [63:0] out_reg_6;
  wire[63:0] T7;
  reg [63:0] out_reg_7;
  wire[63:0] T8;
  reg [63:0] out_reg_8;
  wire[63:0] T9;
  reg [63:0] out_reg_9;
  wire[63:0] T10;
  reg [63:0] out_reg_10;
  wire[63:0] T11;
  reg [63:0] out_reg_11;
  wire[63:0] T12;
  reg [63:0] out_reg_12;
  wire[63:0] T13;
  reg [63:0] out_reg_13;
  wire[63:0] T14;
  reg [63:0] out_reg_14;
  wire[63:0] T15;
  reg [63:0] out_reg_15;
  wire[63:0] T16;
  reg  start_next_stage_reg;
  wire T19;
  wire T17;
  wire T18;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    out_reg_0 = {2{$random}};
    out_reg_1 = {2{$random}};
    out_reg_2 = {2{$random}};
    out_reg_3 = {2{$random}};
    out_reg_4 = {2{$random}};
    out_reg_5 = {2{$random}};
    out_reg_6 = {2{$random}};
    out_reg_7 = {2{$random}};
    out_reg_8 = {2{$random}};
    out_reg_9 = {2{$random}};
    out_reg_10 = {2{$random}};
    out_reg_11 = {2{$random}};
    out_reg_12 = {2{$random}};
    out_reg_13 = {2{$random}};
    out_reg_14 = {2{$random}};
    out_reg_15 = {2{$random}};
    start_next_stage_reg = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_out_0 = out_reg_0;
  assign T0 = T1 ? io_in_0 : out_reg_0;
  assign T1 = io_clk_en & io_start;
  assign io_out_1 = out_reg_1;
  assign T2 = T1 ? io_in_8 : out_reg_1;
  assign io_out_2 = out_reg_2;
  assign T3 = T1 ? io_in_2 : out_reg_2;
  assign io_out_3 = out_reg_3;
  assign T4 = T1 ? io_in_10 : out_reg_3;
  assign io_out_4 = out_reg_4;
  assign T5 = T1 ? io_in_4 : out_reg_4;
  assign io_out_5 = out_reg_5;
  assign T6 = T1 ? io_in_12 : out_reg_5;
  assign io_out_6 = out_reg_6;
  assign T7 = T1 ? io_in_6 : out_reg_6;
  assign io_out_7 = out_reg_7;
  assign T8 = T1 ? io_in_14 : out_reg_7;
  assign io_out_8 = out_reg_8;
  assign T9 = T1 ? io_in_1 : out_reg_8;
  assign io_out_9 = out_reg_9;
  assign T10 = T1 ? io_in_9 : out_reg_9;
  assign io_out_10 = out_reg_10;
  assign T11 = T1 ? io_in_3 : out_reg_10;
  assign io_out_11 = out_reg_11;
  assign T12 = T1 ? io_in_11 : out_reg_11;
  assign io_out_12 = out_reg_12;
  assign T13 = T1 ? io_in_5 : out_reg_12;
  assign io_out_13 = out_reg_13;
  assign T14 = T1 ? io_in_13 : out_reg_13;
  assign io_out_14 = out_reg_14;
  assign T15 = T1 ? io_in_7 : out_reg_14;
  assign io_out_15 = out_reg_15;
  assign T16 = T1 ? io_in_15 : out_reg_15;
  assign io_start_next_stage = start_next_stage_reg;
  assign T19 = reset ? 1'h0 : T17;
  assign T17 = T18 ? 1'h1 : start_next_stage_reg;
  assign T18 = io_start & io_clk_en;

  always @(posedge clk) begin
    if(T1) begin
      out_reg_0 <= io_in_0;
    end
    if(T1) begin
      out_reg_1 <= io_in_8;
    end
    if(T1) begin
      out_reg_2 <= io_in_2;
    end
    if(T1) begin
      out_reg_3 <= io_in_10;
    end
    if(T1) begin
      out_reg_4 <= io_in_4;
    end
    if(T1) begin
      out_reg_5 <= io_in_12;
    end
    if(T1) begin
      out_reg_6 <= io_in_6;
    end
    if(T1) begin
      out_reg_7 <= io_in_14;
    end
    if(T1) begin
      out_reg_8 <= io_in_1;
    end
    if(T1) begin
      out_reg_9 <= io_in_9;
    end
    if(T1) begin
      out_reg_10 <= io_in_3;
    end
    if(T1) begin
      out_reg_11 <= io_in_11;
    end
    if(T1) begin
      out_reg_12 <= io_in_5;
    end
    if(T1) begin
      out_reg_13 <= io_in_13;
    end
    if(T1) begin
      out_reg_14 <= io_in_7;
    end
    if(T1) begin
      out_reg_15 <= io_in_15;
    end
    if(reset) begin
      start_next_stage_reg <= 1'h0;
    end else if(T18) begin
      start_next_stage_reg <= 1'h1;
    end
  end
endmodule

module crossbarShiftDown(input clk, input reset,
    input  io_clk_en,
    input  io_start,
    output io_start_next_stage,
    input [63:0] io_in_15,
    input [63:0] io_in_14,
    input [63:0] io_in_13,
    input [63:0] io_in_12,
    input [63:0] io_in_11,
    input [63:0] io_in_10,
    input [63:0] io_in_9,
    input [63:0] io_in_8,
    input [63:0] io_in_7,
    input [63:0] io_in_6,
    input [63:0] io_in_5,
    input [63:0] io_in_4,
    input [63:0] io_in_3,
    input [63:0] io_in_2,
    input [63:0] io_in_1,
    input [63:0] io_in_0,
    output[63:0] io_out_15,
    output[63:0] io_out_14,
    output[63:0] io_out_13,
    output[63:0] io_out_12,
    output[63:0] io_out_11,
    output[63:0] io_out_10,
    output[63:0] io_out_9,
    output[63:0] io_out_8,
    output[63:0] io_out_7,
    output[63:0] io_out_6,
    output[63:0] io_out_5,
    output[63:0] io_out_4,
    output[63:0] io_out_3,
    output[63:0] io_out_2,
    output[63:0] io_out_1,
    output[63:0] io_out_0
);

  reg [63:0] out_reg_0;
  wire[63:0] T0;
  wire[63:0] T1;
  wire[63:0] T2;
  wire[63:0] T3;
  wire T4;
  wire T5;
  reg [1:0] timestamp;
  wire[1:0] T77;
  wire[1:0] T6;
  wire[1:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  reg [63:0] out_reg_1;
  wire[63:0] T16;
  wire[63:0] T17;
  wire[63:0] T18;
  wire[63:0] T19;
  reg [63:0] out_reg_2;
  wire[63:0] T20;
  wire[63:0] T21;
  wire[63:0] T22;
  wire[63:0] T23;
  reg [63:0] out_reg_3;
  wire[63:0] T24;
  wire[63:0] T25;
  wire[63:0] T26;
  wire[63:0] T27;
  reg [63:0] out_reg_4;
  wire[63:0] T28;
  wire[63:0] T29;
  wire[63:0] T30;
  wire[63:0] T31;
  reg [63:0] out_reg_5;
  wire[63:0] T32;
  wire[63:0] T33;
  wire[63:0] T34;
  wire[63:0] T35;
  reg [63:0] out_reg_6;
  wire[63:0] T36;
  wire[63:0] T37;
  wire[63:0] T38;
  wire[63:0] T39;
  reg [63:0] out_reg_7;
  wire[63:0] T40;
  wire[63:0] T41;
  wire[63:0] T42;
  wire[63:0] T43;
  reg [63:0] out_reg_8;
  wire[63:0] T44;
  wire[63:0] T45;
  wire[63:0] T46;
  wire[63:0] T47;
  reg [63:0] out_reg_9;
  wire[63:0] T48;
  wire[63:0] T49;
  wire[63:0] T50;
  wire[63:0] T51;
  reg [63:0] out_reg_10;
  wire[63:0] T52;
  wire[63:0] T53;
  wire[63:0] T54;
  wire[63:0] T55;
  reg [63:0] out_reg_11;
  wire[63:0] T56;
  wire[63:0] T57;
  wire[63:0] T58;
  wire[63:0] T59;
  reg [63:0] out_reg_12;
  wire[63:0] T60;
  wire[63:0] T61;
  wire[63:0] T62;
  wire[63:0] T63;
  reg [63:0] out_reg_13;
  wire[63:0] T64;
  wire[63:0] T65;
  wire[63:0] T66;
  wire[63:0] T67;
  reg [63:0] out_reg_14;
  wire[63:0] T68;
  wire[63:0] T69;
  wire[63:0] T70;
  wire[63:0] T71;
  reg [63:0] out_reg_15;
  wire[63:0] T72;
  wire[63:0] T73;
  wire[63:0] T74;
  wire[63:0] T75;
  reg  start_next_stage_reg;
  wire T78;
  wire T76;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    out_reg_0 = {2{$random}};
    timestamp = {1{$random}};
    out_reg_1 = {2{$random}};
    out_reg_2 = {2{$random}};
    out_reg_3 = {2{$random}};
    out_reg_4 = {2{$random}};
    out_reg_5 = {2{$random}};
    out_reg_6 = {2{$random}};
    out_reg_7 = {2{$random}};
    out_reg_8 = {2{$random}};
    out_reg_9 = {2{$random}};
    out_reg_10 = {2{$random}};
    out_reg_11 = {2{$random}};
    out_reg_12 = {2{$random}};
    out_reg_13 = {2{$random}};
    out_reg_14 = {2{$random}};
    out_reg_15 = {2{$random}};
    start_next_stage_reg = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_out_0 = out_reg_0;
  assign T0 = T14 ? io_in_10 : T1;
  assign T1 = T12 ? io_in_12 : T2;
  assign T2 = T10 ? io_in_14 : T3;
  assign T3 = T4 ? io_in_0 : out_reg_0;
  assign T4 = T9 & T5;
  assign T5 = timestamp == 2'h0;
  assign T77 = reset ? 2'h0 : T6;
  assign T6 = T8 ? T7 : timestamp;
  assign T7 = timestamp + 2'h1;
  assign T8 = io_clk_en & io_start;
  assign T9 = io_start & io_clk_en;
  assign T10 = T9 & T11;
  assign T11 = timestamp == 2'h1;
  assign T12 = T9 & T13;
  assign T13 = timestamp == 2'h2;
  assign T14 = T9 & T15;
  assign T15 = timestamp == 2'h3;
  assign io_out_1 = out_reg_1;
  assign T16 = T14 ? io_in_11 : T17;
  assign T17 = T12 ? io_in_13 : T18;
  assign T18 = T10 ? io_in_15 : T19;
  assign T19 = T4 ? io_in_1 : out_reg_1;
  assign io_out_2 = out_reg_2;
  assign T20 = T14 ? io_in_12 : T21;
  assign T21 = T12 ? io_in_14 : T22;
  assign T22 = T10 ? io_in_0 : T23;
  assign T23 = T4 ? io_in_2 : out_reg_2;
  assign io_out_3 = out_reg_3;
  assign T24 = T14 ? io_in_13 : T25;
  assign T25 = T12 ? io_in_15 : T26;
  assign T26 = T10 ? io_in_1 : T27;
  assign T27 = T4 ? io_in_3 : out_reg_3;
  assign io_out_4 = out_reg_4;
  assign T28 = T14 ? io_in_14 : T29;
  assign T29 = T12 ? io_in_0 : T30;
  assign T30 = T10 ? io_in_2 : T31;
  assign T31 = T4 ? io_in_4 : out_reg_4;
  assign io_out_5 = out_reg_5;
  assign T32 = T14 ? io_in_15 : T33;
  assign T33 = T12 ? io_in_1 : T34;
  assign T34 = T10 ? io_in_3 : T35;
  assign T35 = T4 ? io_in_5 : out_reg_5;
  assign io_out_6 = out_reg_6;
  assign T36 = T14 ? io_in_0 : T37;
  assign T37 = T12 ? io_in_2 : T38;
  assign T38 = T10 ? io_in_4 : T39;
  assign T39 = T4 ? io_in_6 : out_reg_6;
  assign io_out_7 = out_reg_7;
  assign T40 = T14 ? io_in_1 : T41;
  assign T41 = T12 ? io_in_3 : T42;
  assign T42 = T10 ? io_in_5 : T43;
  assign T43 = T4 ? io_in_7 : out_reg_7;
  assign io_out_8 = out_reg_8;
  assign T44 = T14 ? io_in_2 : T45;
  assign T45 = T12 ? io_in_4 : T46;
  assign T46 = T10 ? io_in_6 : T47;
  assign T47 = T4 ? io_in_8 : out_reg_8;
  assign io_out_9 = out_reg_9;
  assign T48 = T14 ? io_in_3 : T49;
  assign T49 = T12 ? io_in_5 : T50;
  assign T50 = T10 ? io_in_7 : T51;
  assign T51 = T4 ? io_in_9 : out_reg_9;
  assign io_out_10 = out_reg_10;
  assign T52 = T14 ? io_in_4 : T53;
  assign T53 = T12 ? io_in_6 : T54;
  assign T54 = T10 ? io_in_8 : T55;
  assign T55 = T4 ? io_in_10 : out_reg_10;
  assign io_out_11 = out_reg_11;
  assign T56 = T14 ? io_in_5 : T57;
  assign T57 = T12 ? io_in_7 : T58;
  assign T58 = T10 ? io_in_9 : T59;
  assign T59 = T4 ? io_in_11 : out_reg_11;
  assign io_out_12 = out_reg_12;
  assign T60 = T14 ? io_in_6 : T61;
  assign T61 = T12 ? io_in_8 : T62;
  assign T62 = T10 ? io_in_10 : T63;
  assign T63 = T4 ? io_in_12 : out_reg_12;
  assign io_out_13 = out_reg_13;
  assign T64 = T14 ? io_in_7 : T65;
  assign T65 = T12 ? io_in_9 : T66;
  assign T66 = T10 ? io_in_11 : T67;
  assign T67 = T4 ? io_in_13 : out_reg_13;
  assign io_out_14 = out_reg_14;
  assign T68 = T14 ? io_in_8 : T69;
  assign T69 = T12 ? io_in_10 : T70;
  assign T70 = T10 ? io_in_12 : T71;
  assign T71 = T4 ? io_in_14 : out_reg_14;
  assign io_out_15 = out_reg_15;
  assign T72 = T14 ? io_in_9 : T73;
  assign T73 = T12 ? io_in_11 : T74;
  assign T74 = T10 ? io_in_13 : T75;
  assign T75 = T4 ? io_in_15 : out_reg_15;
  assign io_start_next_stage = start_next_stage_reg;
  assign T78 = reset ? 1'h0 : T76;
  assign T76 = T8 ? 1'h1 : start_next_stage_reg;

  always @(posedge clk) begin
    if(T14) begin
      out_reg_0 <= io_in_10;
    end else if(T12) begin
      out_reg_0 <= io_in_12;
    end else if(T10) begin
      out_reg_0 <= io_in_14;
    end else if(T4) begin
      out_reg_0 <= io_in_0;
    end
    if(reset) begin
      timestamp <= 2'h0;
    end else if(T8) begin
      timestamp <= T7;
    end
    if(T14) begin
      out_reg_1 <= io_in_11;
    end else if(T12) begin
      out_reg_1 <= io_in_13;
    end else if(T10) begin
      out_reg_1 <= io_in_15;
    end else if(T4) begin
      out_reg_1 <= io_in_1;
    end
    if(T14) begin
      out_reg_2 <= io_in_12;
    end else if(T12) begin
      out_reg_2 <= io_in_14;
    end else if(T10) begin
      out_reg_2 <= io_in_0;
    end else if(T4) begin
      out_reg_2 <= io_in_2;
    end
    if(T14) begin
      out_reg_3 <= io_in_13;
    end else if(T12) begin
      out_reg_3 <= io_in_15;
    end else if(T10) begin
      out_reg_3 <= io_in_1;
    end else if(T4) begin
      out_reg_3 <= io_in_3;
    end
    if(T14) begin
      out_reg_4 <= io_in_14;
    end else if(T12) begin
      out_reg_4 <= io_in_0;
    end else if(T10) begin
      out_reg_4 <= io_in_2;
    end else if(T4) begin
      out_reg_4 <= io_in_4;
    end
    if(T14) begin
      out_reg_5 <= io_in_15;
    end else if(T12) begin
      out_reg_5 <= io_in_1;
    end else if(T10) begin
      out_reg_5 <= io_in_3;
    end else if(T4) begin
      out_reg_5 <= io_in_5;
    end
    if(T14) begin
      out_reg_6 <= io_in_0;
    end else if(T12) begin
      out_reg_6 <= io_in_2;
    end else if(T10) begin
      out_reg_6 <= io_in_4;
    end else if(T4) begin
      out_reg_6 <= io_in_6;
    end
    if(T14) begin
      out_reg_7 <= io_in_1;
    end else if(T12) begin
      out_reg_7 <= io_in_3;
    end else if(T10) begin
      out_reg_7 <= io_in_5;
    end else if(T4) begin
      out_reg_7 <= io_in_7;
    end
    if(T14) begin
      out_reg_8 <= io_in_2;
    end else if(T12) begin
      out_reg_8 <= io_in_4;
    end else if(T10) begin
      out_reg_8 <= io_in_6;
    end else if(T4) begin
      out_reg_8 <= io_in_8;
    end
    if(T14) begin
      out_reg_9 <= io_in_3;
    end else if(T12) begin
      out_reg_9 <= io_in_5;
    end else if(T10) begin
      out_reg_9 <= io_in_7;
    end else if(T4) begin
      out_reg_9 <= io_in_9;
    end
    if(T14) begin
      out_reg_10 <= io_in_4;
    end else if(T12) begin
      out_reg_10 <= io_in_6;
    end else if(T10) begin
      out_reg_10 <= io_in_8;
    end else if(T4) begin
      out_reg_10 <= io_in_10;
    end
    if(T14) begin
      out_reg_11 <= io_in_5;
    end else if(T12) begin
      out_reg_11 <= io_in_7;
    end else if(T10) begin
      out_reg_11 <= io_in_9;
    end else if(T4) begin
      out_reg_11 <= io_in_11;
    end
    if(T14) begin
      out_reg_12 <= io_in_6;
    end else if(T12) begin
      out_reg_12 <= io_in_8;
    end else if(T10) begin
      out_reg_12 <= io_in_10;
    end else if(T4) begin
      out_reg_12 <= io_in_12;
    end
    if(T14) begin
      out_reg_13 <= io_in_7;
    end else if(T12) begin
      out_reg_13 <= io_in_9;
    end else if(T10) begin
      out_reg_13 <= io_in_11;
    end else if(T4) begin
      out_reg_13 <= io_in_13;
    end
    if(T14) begin
      out_reg_14 <= io_in_8;
    end else if(T12) begin
      out_reg_14 <= io_in_10;
    end else if(T10) begin
      out_reg_14 <= io_in_12;
    end else if(T4) begin
      out_reg_14 <= io_in_14;
    end
    if(T14) begin
      out_reg_15 <= io_in_9;
    end else if(T12) begin
      out_reg_15 <= io_in_11;
    end else if(T10) begin
      out_reg_15 <= io_in_13;
    end else if(T4) begin
      out_reg_15 <= io_in_15;
    end
    if(reset) begin
      start_next_stage_reg <= 1'h0;
    end else if(T8) begin
      start_next_stage_reg <= 1'h1;
    end
  end
endmodule

module single_port_ram(input clk,
    input [63:0] io_data,
    input [1:0] io_addr,
    input  io_we,
    output[63:0] io_q
);

  reg [63:0] out;
  wire[63:0] T0;
  wire[63:0] T1;
  reg [63:0] myMem [3:0];
  wire[63:0] T2;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    out = {2{$random}};
    for (initvar = 0; initvar < 4; initvar = initvar+1)
      myMem[initvar] = {2{$random}};
  end
// synthesis translate_on
`endif

  assign io_q = out;
  assign T0 = io_we ? T1 : out;
  assign T1 = myMem[io_addr];

  always @(posedge clk) begin
    if(io_we) begin
      out <= T1;
    end
    if (io_we)
      myMem[io_addr] <= io_data;
  end
endmodule

module memArray(input clk, input reset,
    input  io_clk_en,
    input  io_start,
    output io_start_next_stage,
    input [63:0] io_in_15,
    input [63:0] io_in_14,
    input [63:0] io_in_13,
    input [63:0] io_in_12,
    input [63:0] io_in_11,
    input [63:0] io_in_10,
    input [63:0] io_in_9,
    input [63:0] io_in_8,
    input [63:0] io_in_7,
    input [63:0] io_in_6,
    input [63:0] io_in_5,
    input [63:0] io_in_4,
    input [63:0] io_in_3,
    input [63:0] io_in_2,
    input [63:0] io_in_1,
    input [63:0] io_in_0,
    output[63:0] io_out_15,
    output[63:0] io_out_14,
    output[63:0] io_out_13,
    output[63:0] io_out_12,
    output[63:0] io_out_11,
    output[63:0] io_out_10,
    output[63:0] io_out_9,
    output[63:0] io_out_8,
    output[63:0] io_out_7,
    output[63:0] io_out_6,
    output[63:0] io_out_5,
    output[63:0] io_out_4,
    output[63:0] io_out_3,
    output[63:0] io_out_2,
    output[63:0] io_out_1,
    output[63:0] io_out_0
);

  wire T0;
  reg [1:0] address_7;
  wire[1:0] T105;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire[1:0] T6;
  wire T7;
  wire T8;
  reg [1:0] state;
  wire[1:0] T106;
  wire[1:0] T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire T14;
  reg [1:0] counter;
  wire[1:0] T107;
  wire[1:0] T15;
  wire[1:0] T16;
  wire[1:0] T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire[1:0] T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[1:0] T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire[1:0] T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  reg [1:0] address_6;
  wire[1:0] T108;
  wire[1:0] T35;
  wire[1:0] T36;
  wire[1:0] T37;
  wire[1:0] T38;
  wire[1:0] T39;
  wire[1:0] T40;
  wire[1:0] T41;
  wire[1:0] T42;
  wire T43;
  wire T44;
  reg [1:0] address_5;
  wire[1:0] T109;
  wire[1:0] T45;
  wire[1:0] T46;
  wire[1:0] T47;
  wire[1:0] T48;
  wire[1:0] T49;
  wire[1:0] T50;
  wire[1:0] T51;
  wire[1:0] T52;
  wire T53;
  wire T54;
  reg [1:0] address_4;
  wire[1:0] T110;
  wire[1:0] T55;
  wire[1:0] T56;
  wire[1:0] T57;
  wire[1:0] T58;
  wire[1:0] T59;
  wire[1:0] T60;
  wire[1:0] T61;
  wire[1:0] T62;
  wire T63;
  wire T64;
  reg [1:0] address_3;
  wire[1:0] T111;
  wire[1:0] T65;
  wire[1:0] T66;
  wire[1:0] T67;
  wire[1:0] T68;
  wire[1:0] T69;
  wire[1:0] T70;
  wire[1:0] T71;
  wire[1:0] T72;
  wire T73;
  wire T74;
  reg [1:0] address_2;
  wire[1:0] T112;
  wire[1:0] T75;
  wire[1:0] T76;
  wire[1:0] T77;
  wire[1:0] T78;
  wire[1:0] T79;
  wire[1:0] T80;
  wire[1:0] T81;
  wire[1:0] T82;
  wire T83;
  wire T84;
  reg [1:0] address_1;
  wire[1:0] T113;
  wire[1:0] T85;
  wire[1:0] T86;
  wire[1:0] T87;
  wire[1:0] T88;
  wire[1:0] T89;
  wire[1:0] T90;
  wire[1:0] T91;
  wire[1:0] T92;
  wire T93;
  wire T94;
  reg [1:0] address_0;
  wire[1:0] T114;
  wire[1:0] T95;
  wire[1:0] T96;
  wire[1:0] T97;
  wire[1:0] T98;
  wire[1:0] T99;
  wire[1:0] T100;
  wire[1:0] T101;
  wire[1:0] T102;
  wire T103;
  reg  start_next_stage_reg;
  wire T115;
  wire T104;
  wire[63:0] single_port_ram_io_q;
  wire[63:0] single_port_ram_1_io_q;
  wire[63:0] single_port_ram_2_io_q;
  wire[63:0] single_port_ram_3_io_q;
  wire[63:0] single_port_ram_4_io_q;
  wire[63:0] single_port_ram_5_io_q;
  wire[63:0] single_port_ram_6_io_q;
  wire[63:0] single_port_ram_7_io_q;
  wire[63:0] single_port_ram_8_io_q;
  wire[63:0] single_port_ram_9_io_q;
  wire[63:0] single_port_ram_10_io_q;
  wire[63:0] single_port_ram_11_io_q;
  wire[63:0] single_port_ram_12_io_q;
  wire[63:0] single_port_ram_13_io_q;
  wire[63:0] single_port_ram_14_io_q;
  wire[63:0] single_port_ram_15_io_q;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    address_7 = {1{$random}};
    state = {1{$random}};
    counter = {1{$random}};
    address_6 = {1{$random}};
    address_5 = {1{$random}};
    address_4 = {1{$random}};
    address_3 = {1{$random}};
    address_2 = {1{$random}};
    address_1 = {1{$random}};
    address_0 = {1{$random}};
    start_next_stage_reg = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_start & io_clk_en;
  assign T105 = reset ? 2'h0 : T1;
  assign T1 = T31 ? T30 : T2;
  assign T2 = T28 ? 2'h0 : T3;
  assign T3 = T26 ? T25 : T4;
  assign T4 = T13 ? 2'h3 : T5;
  assign T5 = T7 ? T6 : address_7;
  assign T6 = address_7 + 2'h1;
  assign T7 = T12 & T8;
  assign T8 = state == 2'h0;
  assign T106 = reset ? 2'h0 : T9;
  assign T9 = T28 ? 2'h1 : T10;
  assign T10 = T13 ? 2'h2 : T11;
  assign T11 = T7 ? 2'h1 : state;
  assign T12 = io_clk_en & io_start;
  assign T13 = T23 & T14;
  assign T14 = counter == 2'h3;
  assign T107 = reset ? 2'h0 : T15;
  assign T15 = T21 ? T20 : T16;
  assign T16 = T23 ? T19 : T17;
  assign T17 = T7 ? T18 : counter;
  assign T18 = counter + 2'h1;
  assign T19 = counter + 2'h1;
  assign T20 = counter + 2'h1;
  assign T21 = T12 & T22;
  assign T22 = state == 2'h2;
  assign T23 = T12 & T24;
  assign T24 = state == 2'h1;
  assign T25 = address_7 + 2'h1;
  assign T26 = T23 & T27;
  assign T27 = T14 ^ 1'h1;
  assign T28 = T21 & T29;
  assign T29 = counter == 2'h3;
  assign T30 = address_7 - 2'h1;
  assign T31 = T21 & T32;
  assign T32 = T29 ^ 1'h1;
  assign T33 = io_start & io_clk_en;
  assign T34 = io_start & io_clk_en;
  assign T108 = reset ? 2'h0 : T35;
  assign T35 = T31 ? T42 : T36;
  assign T36 = T28 ? 2'h0 : T37;
  assign T37 = T26 ? T41 : T38;
  assign T38 = T13 ? 2'h2 : T39;
  assign T39 = T7 ? T40 : address_6;
  assign T40 = address_6 + 2'h1;
  assign T41 = address_6 + 2'h1;
  assign T42 = address_6 - 2'h1;
  assign T43 = io_start & io_clk_en;
  assign T44 = io_start & io_clk_en;
  assign T109 = reset ? 2'h0 : T45;
  assign T45 = T31 ? T52 : T46;
  assign T46 = T28 ? 2'h0 : T47;
  assign T47 = T26 ? T51 : T48;
  assign T48 = T13 ? 2'h1 : T49;
  assign T49 = T7 ? T50 : address_5;
  assign T50 = address_5 + 2'h1;
  assign T51 = address_5 + 2'h1;
  assign T52 = address_5 - 2'h1;
  assign T53 = io_start & io_clk_en;
  assign T54 = io_start & io_clk_en;
  assign T110 = reset ? 2'h0 : T55;
  assign T55 = T31 ? T62 : T56;
  assign T56 = T28 ? 2'h0 : T57;
  assign T57 = T26 ? T61 : T58;
  assign T58 = T13 ? 2'h0 : T59;
  assign T59 = T7 ? T60 : address_4;
  assign T60 = address_4 + 2'h1;
  assign T61 = address_4 + 2'h1;
  assign T62 = address_4 - 2'h1;
  assign T63 = io_start & io_clk_en;
  assign T64 = io_start & io_clk_en;
  assign T111 = reset ? 2'h0 : T65;
  assign T65 = T31 ? T72 : T66;
  assign T66 = T28 ? 2'h0 : T67;
  assign T67 = T26 ? T71 : T68;
  assign T68 = T13 ? 2'h3 : T69;
  assign T69 = T7 ? T70 : address_3;
  assign T70 = address_3 + 2'h1;
  assign T71 = address_3 + 2'h1;
  assign T72 = address_3 - 2'h1;
  assign T73 = io_start & io_clk_en;
  assign T74 = io_start & io_clk_en;
  assign T112 = reset ? 2'h0 : T75;
  assign T75 = T31 ? T82 : T76;
  assign T76 = T28 ? 2'h0 : T77;
  assign T77 = T26 ? T81 : T78;
  assign T78 = T13 ? 2'h2 : T79;
  assign T79 = T7 ? T80 : address_2;
  assign T80 = address_2 + 2'h1;
  assign T81 = address_2 + 2'h1;
  assign T82 = address_2 - 2'h1;
  assign T83 = io_start & io_clk_en;
  assign T84 = io_start & io_clk_en;
  assign T113 = reset ? 2'h0 : T85;
  assign T85 = T31 ? T92 : T86;
  assign T86 = T28 ? 2'h0 : T87;
  assign T87 = T26 ? T91 : T88;
  assign T88 = T13 ? 2'h1 : T89;
  assign T89 = T7 ? T90 : address_1;
  assign T90 = address_1 + 2'h1;
  assign T91 = address_1 + 2'h1;
  assign T92 = address_1 - 2'h1;
  assign T93 = io_start & io_clk_en;
  assign T94 = io_start & io_clk_en;
  assign T114 = reset ? 2'h0 : T95;
  assign T95 = T31 ? T102 : T96;
  assign T96 = T28 ? 2'h0 : T97;
  assign T97 = T26 ? T101 : T98;
  assign T98 = T13 ? 2'h0 : T99;
  assign T99 = T7 ? T100 : address_0;
  assign T100 = address_0 + 2'h1;
  assign T101 = address_0 + 2'h1;
  assign T102 = address_0 - 2'h1;
  assign T103 = io_start & io_clk_en;
  assign io_out_0 = single_port_ram_io_q;
  assign io_out_1 = single_port_ram_1_io_q;
  assign io_out_2 = single_port_ram_2_io_q;
  assign io_out_3 = single_port_ram_3_io_q;
  assign io_out_4 = single_port_ram_4_io_q;
  assign io_out_5 = single_port_ram_5_io_q;
  assign io_out_6 = single_port_ram_6_io_q;
  assign io_out_7 = single_port_ram_7_io_q;
  assign io_out_8 = single_port_ram_8_io_q;
  assign io_out_9 = single_port_ram_9_io_q;
  assign io_out_10 = single_port_ram_10_io_q;
  assign io_out_11 = single_port_ram_11_io_q;
  assign io_out_12 = single_port_ram_12_io_q;
  assign io_out_13 = single_port_ram_13_io_q;
  assign io_out_14 = single_port_ram_14_io_q;
  assign io_out_15 = single_port_ram_15_io_q;
  assign io_start_next_stage = start_next_stage_reg;
  assign T115 = reset ? 1'h0 : T104;
  assign T104 = T21 ? 1'h1 : start_next_stage_reg;
  single_port_ram single_port_ram(.clk(clk),
       .io_data( io_in_0 ),
       .io_addr( address_0 ),
       .io_we( T103 ),
       .io_q( single_port_ram_io_q )
  );
  single_port_ram single_port_ram_1(.clk(clk),
       .io_data( io_in_1 ),
       .io_addr( address_0 ),
       .io_we( T94 ),
       .io_q( single_port_ram_1_io_q )
  );
  single_port_ram single_port_ram_2(.clk(clk),
       .io_data( io_in_2 ),
       .io_addr( address_1 ),
       .io_we( T93 ),
       .io_q( single_port_ram_2_io_q )
  );
  single_port_ram single_port_ram_3(.clk(clk),
       .io_data( io_in_3 ),
       .io_addr( address_1 ),
       .io_we( T84 ),
       .io_q( single_port_ram_3_io_q )
  );
  single_port_ram single_port_ram_4(.clk(clk),
       .io_data( io_in_4 ),
       .io_addr( address_2 ),
       .io_we( T83 ),
       .io_q( single_port_ram_4_io_q )
  );
  single_port_ram single_port_ram_5(.clk(clk),
       .io_data( io_in_5 ),
       .io_addr( address_2 ),
       .io_we( T74 ),
       .io_q( single_port_ram_5_io_q )
  );
  single_port_ram single_port_ram_6(.clk(clk),
       .io_data( io_in_6 ),
       .io_addr( address_3 ),
       .io_we( T73 ),
       .io_q( single_port_ram_6_io_q )
  );
  single_port_ram single_port_ram_7(.clk(clk),
       .io_data( io_in_7 ),
       .io_addr( address_3 ),
       .io_we( T64 ),
       .io_q( single_port_ram_7_io_q )
  );
  single_port_ram single_port_ram_8(.clk(clk),
       .io_data( io_in_8 ),
       .io_addr( address_4 ),
       .io_we( T63 ),
       .io_q( single_port_ram_8_io_q )
  );
  single_port_ram single_port_ram_9(.clk(clk),
       .io_data( io_in_9 ),
       .io_addr( address_4 ),
       .io_we( T54 ),
       .io_q( single_port_ram_9_io_q )
  );
  single_port_ram single_port_ram_10(.clk(clk),
       .io_data( io_in_10 ),
       .io_addr( address_5 ),
       .io_we( T53 ),
       .io_q( single_port_ram_10_io_q )
  );
  single_port_ram single_port_ram_11(.clk(clk),
       .io_data( io_in_11 ),
       .io_addr( address_5 ),
       .io_we( T44 ),
       .io_q( single_port_ram_11_io_q )
  );
  single_port_ram single_port_ram_12(.clk(clk),
       .io_data( io_in_12 ),
       .io_addr( address_6 ),
       .io_we( T43 ),
       .io_q( single_port_ram_12_io_q )
  );
  single_port_ram single_port_ram_13(.clk(clk),
       .io_data( io_in_13 ),
       .io_addr( address_6 ),
       .io_we( T34 ),
       .io_q( single_port_ram_13_io_q )
  );
  single_port_ram single_port_ram_14(.clk(clk),
       .io_data( io_in_14 ),
       .io_addr( address_7 ),
       .io_we( T33 ),
       .io_q( single_port_ram_14_io_q )
  );
  single_port_ram single_port_ram_15(.clk(clk),
       .io_data( io_in_15 ),
       .io_addr( address_7 ),
       .io_we( T0 ),
       .io_q( single_port_ram_15_io_q )
  );

  always @(posedge clk) begin
    if(reset) begin
      address_7 <= 2'h0;
    end else if(T31) begin
      address_7 <= T30;
    end else if(T28) begin
      address_7 <= 2'h0;
    end else if(T26) begin
      address_7 <= T25;
    end else if(T13) begin
      address_7 <= 2'h3;
    end else if(T7) begin
      address_7 <= T6;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(T28) begin
      state <= 2'h1;
    end else if(T13) begin
      state <= 2'h2;
    end else if(T7) begin
      state <= 2'h1;
    end
    if(reset) begin
      counter <= 2'h0;
    end else if(T21) begin
      counter <= T20;
    end else if(T23) begin
      counter <= T19;
    end else if(T7) begin
      counter <= T18;
    end
    if(reset) begin
      address_6 <= 2'h0;
    end else if(T31) begin
      address_6 <= T42;
    end else if(T28) begin
      address_6 <= 2'h0;
    end else if(T26) begin
      address_6 <= T41;
    end else if(T13) begin
      address_6 <= 2'h2;
    end else if(T7) begin
      address_6 <= T40;
    end
    if(reset) begin
      address_5 <= 2'h0;
    end else if(T31) begin
      address_5 <= T52;
    end else if(T28) begin
      address_5 <= 2'h0;
    end else if(T26) begin
      address_5 <= T51;
    end else if(T13) begin
      address_5 <= 2'h1;
    end else if(T7) begin
      address_5 <= T50;
    end
    if(reset) begin
      address_4 <= 2'h0;
    end else if(T31) begin
      address_4 <= T62;
    end else if(T28) begin
      address_4 <= 2'h0;
    end else if(T26) begin
      address_4 <= T61;
    end else if(T13) begin
      address_4 <= 2'h0;
    end else if(T7) begin
      address_4 <= T60;
    end
    if(reset) begin
      address_3 <= 2'h0;
    end else if(T31) begin
      address_3 <= T72;
    end else if(T28) begin
      address_3 <= 2'h0;
    end else if(T26) begin
      address_3 <= T71;
    end else if(T13) begin
      address_3 <= 2'h3;
    end else if(T7) begin
      address_3 <= T70;
    end
    if(reset) begin
      address_2 <= 2'h0;
    end else if(T31) begin
      address_2 <= T82;
    end else if(T28) begin
      address_2 <= 2'h0;
    end else if(T26) begin
      address_2 <= T81;
    end else if(T13) begin
      address_2 <= 2'h2;
    end else if(T7) begin
      address_2 <= T80;
    end
    if(reset) begin
      address_1 <= 2'h0;
    end else if(T31) begin
      address_1 <= T92;
    end else if(T28) begin
      address_1 <= 2'h0;
    end else if(T26) begin
      address_1 <= T91;
    end else if(T13) begin
      address_1 <= 2'h1;
    end else if(T7) begin
      address_1 <= T90;
    end
    if(reset) begin
      address_0 <= 2'h0;
    end else if(T31) begin
      address_0 <= T102;
    end else if(T28) begin
      address_0 <= 2'h0;
    end else if(T26) begin
      address_0 <= T101;
    end else if(T13) begin
      address_0 <= 2'h0;
    end else if(T7) begin
      address_0 <= T100;
    end
    if(reset) begin
      start_next_stage_reg <= 1'h0;
    end else if(T21) begin
      start_next_stage_reg <= 1'h1;
    end
  end
endmodule

module crossbarShiftUp(input clk, input reset,
    input  io_clk_en,
    input  io_start,
    output io_start_next_stage,
    input [63:0] io_in_15,
    input [63:0] io_in_14,
    input [63:0] io_in_13,
    input [63:0] io_in_12,
    input [63:0] io_in_11,
    input [63:0] io_in_10,
    input [63:0] io_in_9,
    input [63:0] io_in_8,
    input [63:0] io_in_7,
    input [63:0] io_in_6,
    input [63:0] io_in_5,
    input [63:0] io_in_4,
    input [63:0] io_in_3,
    input [63:0] io_in_2,
    input [63:0] io_in_1,
    input [63:0] io_in_0,
    output[63:0] io_out_15,
    output[63:0] io_out_14,
    output[63:0] io_out_13,
    output[63:0] io_out_12,
    output[63:0] io_out_11,
    output[63:0] io_out_10,
    output[63:0] io_out_9,
    output[63:0] io_out_8,
    output[63:0] io_out_7,
    output[63:0] io_out_6,
    output[63:0] io_out_5,
    output[63:0] io_out_4,
    output[63:0] io_out_3,
    output[63:0] io_out_2,
    output[63:0] io_out_1,
    output[63:0] io_out_0
);

  reg [63:0] out_reg_0;
  wire[63:0] T0;
  wire[63:0] T1;
  wire[63:0] T2;
  wire[63:0] T3;
  wire T4;
  wire T5;
  reg [1:0] timestamp;
  wire[1:0] T77;
  wire[1:0] T6;
  wire[1:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  reg [63:0] out_reg_1;
  wire[63:0] T16;
  wire[63:0] T17;
  wire[63:0] T18;
  wire[63:0] T19;
  reg [63:0] out_reg_2;
  wire[63:0] T20;
  wire[63:0] T21;
  wire[63:0] T22;
  wire[63:0] T23;
  reg [63:0] out_reg_3;
  wire[63:0] T24;
  wire[63:0] T25;
  wire[63:0] T26;
  wire[63:0] T27;
  reg [63:0] out_reg_4;
  wire[63:0] T28;
  wire[63:0] T29;
  wire[63:0] T30;
  wire[63:0] T31;
  reg [63:0] out_reg_5;
  wire[63:0] T32;
  wire[63:0] T33;
  wire[63:0] T34;
  wire[63:0] T35;
  reg [63:0] out_reg_6;
  wire[63:0] T36;
  wire[63:0] T37;
  wire[63:0] T38;
  wire[63:0] T39;
  reg [63:0] out_reg_7;
  wire[63:0] T40;
  wire[63:0] T41;
  wire[63:0] T42;
  wire[63:0] T43;
  reg [63:0] out_reg_8;
  wire[63:0] T44;
  wire[63:0] T45;
  wire[63:0] T46;
  wire[63:0] T47;
  reg [63:0] out_reg_9;
  wire[63:0] T48;
  wire[63:0] T49;
  wire[63:0] T50;
  wire[63:0] T51;
  reg [63:0] out_reg_10;
  wire[63:0] T52;
  wire[63:0] T53;
  wire[63:0] T54;
  wire[63:0] T55;
  reg [63:0] out_reg_11;
  wire[63:0] T56;
  wire[63:0] T57;
  wire[63:0] T58;
  wire[63:0] T59;
  reg [63:0] out_reg_12;
  wire[63:0] T60;
  wire[63:0] T61;
  wire[63:0] T62;
  wire[63:0] T63;
  reg [63:0] out_reg_13;
  wire[63:0] T64;
  wire[63:0] T65;
  wire[63:0] T66;
  wire[63:0] T67;
  reg [63:0] out_reg_14;
  wire[63:0] T68;
  wire[63:0] T69;
  wire[63:0] T70;
  wire[63:0] T71;
  reg [63:0] out_reg_15;
  wire[63:0] T72;
  wire[63:0] T73;
  wire[63:0] T74;
  wire[63:0] T75;
  reg  start_next_stage_reg;
  wire T78;
  wire T76;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    out_reg_0 = {2{$random}};
    timestamp = {1{$random}};
    out_reg_1 = {2{$random}};
    out_reg_2 = {2{$random}};
    out_reg_3 = {2{$random}};
    out_reg_4 = {2{$random}};
    out_reg_5 = {2{$random}};
    out_reg_6 = {2{$random}};
    out_reg_7 = {2{$random}};
    out_reg_8 = {2{$random}};
    out_reg_9 = {2{$random}};
    out_reg_10 = {2{$random}};
    out_reg_11 = {2{$random}};
    out_reg_12 = {2{$random}};
    out_reg_13 = {2{$random}};
    out_reg_14 = {2{$random}};
    out_reg_15 = {2{$random}};
    start_next_stage_reg = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_out_0 = out_reg_0;
  assign T0 = T14 ? io_in_6 : T1;
  assign T1 = T12 ? io_in_4 : T2;
  assign T2 = T10 ? io_in_2 : T3;
  assign T3 = T4 ? io_in_0 : out_reg_0;
  assign T4 = T9 & T5;
  assign T5 = timestamp == 2'h0;
  assign T77 = reset ? 2'h0 : T6;
  assign T6 = T8 ? T7 : timestamp;
  assign T7 = timestamp + 2'h1;
  assign T8 = io_clk_en & io_start;
  assign T9 = io_start & io_clk_en;
  assign T10 = T9 & T11;
  assign T11 = timestamp == 2'h1;
  assign T12 = T9 & T13;
  assign T13 = timestamp == 2'h2;
  assign T14 = T9 & T15;
  assign T15 = timestamp == 2'h3;
  assign io_out_1 = out_reg_1;
  assign T16 = T14 ? io_in_7 : T17;
  assign T17 = T12 ? io_in_5 : T18;
  assign T18 = T10 ? io_in_3 : T19;
  assign T19 = T4 ? io_in_1 : out_reg_1;
  assign io_out_2 = out_reg_2;
  assign T20 = T14 ? io_in_8 : T21;
  assign T21 = T12 ? io_in_6 : T22;
  assign T22 = T10 ? io_in_4 : T23;
  assign T23 = T4 ? io_in_2 : out_reg_2;
  assign io_out_3 = out_reg_3;
  assign T24 = T14 ? io_in_9 : T25;
  assign T25 = T12 ? io_in_7 : T26;
  assign T26 = T10 ? io_in_5 : T27;
  assign T27 = T4 ? io_in_3 : out_reg_3;
  assign io_out_4 = out_reg_4;
  assign T28 = T14 ? io_in_10 : T29;
  assign T29 = T12 ? io_in_8 : T30;
  assign T30 = T10 ? io_in_6 : T31;
  assign T31 = T4 ? io_in_4 : out_reg_4;
  assign io_out_5 = out_reg_5;
  assign T32 = T14 ? io_in_11 : T33;
  assign T33 = T12 ? io_in_9 : T34;
  assign T34 = T10 ? io_in_7 : T35;
  assign T35 = T4 ? io_in_5 : out_reg_5;
  assign io_out_6 = out_reg_6;
  assign T36 = T14 ? io_in_12 : T37;
  assign T37 = T12 ? io_in_10 : T38;
  assign T38 = T10 ? io_in_8 : T39;
  assign T39 = T4 ? io_in_6 : out_reg_6;
  assign io_out_7 = out_reg_7;
  assign T40 = T14 ? io_in_13 : T41;
  assign T41 = T12 ? io_in_11 : T42;
  assign T42 = T10 ? io_in_9 : T43;
  assign T43 = T4 ? io_in_7 : out_reg_7;
  assign io_out_8 = out_reg_8;
  assign T44 = T14 ? io_in_14 : T45;
  assign T45 = T12 ? io_in_12 : T46;
  assign T46 = T10 ? io_in_10 : T47;
  assign T47 = T4 ? io_in_8 : out_reg_8;
  assign io_out_9 = out_reg_9;
  assign T48 = T14 ? io_in_15 : T49;
  assign T49 = T12 ? io_in_13 : T50;
  assign T50 = T10 ? io_in_11 : T51;
  assign T51 = T4 ? io_in_9 : out_reg_9;
  assign io_out_10 = out_reg_10;
  assign T52 = T14 ? io_in_0 : T53;
  assign T53 = T12 ? io_in_14 : T54;
  assign T54 = T10 ? io_in_12 : T55;
  assign T55 = T4 ? io_in_10 : out_reg_10;
  assign io_out_11 = out_reg_11;
  assign T56 = T14 ? io_in_1 : T57;
  assign T57 = T12 ? io_in_15 : T58;
  assign T58 = T10 ? io_in_13 : T59;
  assign T59 = T4 ? io_in_11 : out_reg_11;
  assign io_out_12 = out_reg_12;
  assign T60 = T14 ? io_in_2 : T61;
  assign T61 = T12 ? io_in_0 : T62;
  assign T62 = T10 ? io_in_14 : T63;
  assign T63 = T4 ? io_in_12 : out_reg_12;
  assign io_out_13 = out_reg_13;
  assign T64 = T14 ? io_in_3 : T65;
  assign T65 = T12 ? io_in_1 : T66;
  assign T66 = T10 ? io_in_15 : T67;
  assign T67 = T4 ? io_in_13 : out_reg_13;
  assign io_out_14 = out_reg_14;
  assign T68 = T14 ? io_in_4 : T69;
  assign T69 = T12 ? io_in_2 : T70;
  assign T70 = T10 ? io_in_0 : T71;
  assign T71 = T4 ? io_in_14 : out_reg_14;
  assign io_out_15 = out_reg_15;
  assign T72 = T14 ? io_in_5 : T73;
  assign T73 = T12 ? io_in_3 : T74;
  assign T74 = T10 ? io_in_1 : T75;
  assign T75 = T4 ? io_in_15 : out_reg_15;
  assign io_start_next_stage = start_next_stage_reg;
  assign T78 = reset ? 1'h0 : T76;
  assign T76 = T8 ? 1'h1 : start_next_stage_reg;

  always @(posedge clk) begin
    if(T14) begin
      out_reg_0 <= io_in_6;
    end else if(T12) begin
      out_reg_0 <= io_in_4;
    end else if(T10) begin
      out_reg_0 <= io_in_2;
    end else if(T4) begin
      out_reg_0 <= io_in_0;
    end
    if(reset) begin
      timestamp <= 2'h0;
    end else if(T8) begin
      timestamp <= T7;
    end
    if(T14) begin
      out_reg_1 <= io_in_7;
    end else if(T12) begin
      out_reg_1 <= io_in_5;
    end else if(T10) begin
      out_reg_1 <= io_in_3;
    end else if(T4) begin
      out_reg_1 <= io_in_1;
    end
    if(T14) begin
      out_reg_2 <= io_in_8;
    end else if(T12) begin
      out_reg_2 <= io_in_6;
    end else if(T10) begin
      out_reg_2 <= io_in_4;
    end else if(T4) begin
      out_reg_2 <= io_in_2;
    end
    if(T14) begin
      out_reg_3 <= io_in_9;
    end else if(T12) begin
      out_reg_3 <= io_in_7;
    end else if(T10) begin
      out_reg_3 <= io_in_5;
    end else if(T4) begin
      out_reg_3 <= io_in_3;
    end
    if(T14) begin
      out_reg_4 <= io_in_10;
    end else if(T12) begin
      out_reg_4 <= io_in_8;
    end else if(T10) begin
      out_reg_4 <= io_in_6;
    end else if(T4) begin
      out_reg_4 <= io_in_4;
    end
    if(T14) begin
      out_reg_5 <= io_in_11;
    end else if(T12) begin
      out_reg_5 <= io_in_9;
    end else if(T10) begin
      out_reg_5 <= io_in_7;
    end else if(T4) begin
      out_reg_5 <= io_in_5;
    end
    if(T14) begin
      out_reg_6 <= io_in_12;
    end else if(T12) begin
      out_reg_6 <= io_in_10;
    end else if(T10) begin
      out_reg_6 <= io_in_8;
    end else if(T4) begin
      out_reg_6 <= io_in_6;
    end
    if(T14) begin
      out_reg_7 <= io_in_13;
    end else if(T12) begin
      out_reg_7 <= io_in_11;
    end else if(T10) begin
      out_reg_7 <= io_in_9;
    end else if(T4) begin
      out_reg_7 <= io_in_7;
    end
    if(T14) begin
      out_reg_8 <= io_in_14;
    end else if(T12) begin
      out_reg_8 <= io_in_12;
    end else if(T10) begin
      out_reg_8 <= io_in_10;
    end else if(T4) begin
      out_reg_8 <= io_in_8;
    end
    if(T14) begin
      out_reg_9 <= io_in_15;
    end else if(T12) begin
      out_reg_9 <= io_in_13;
    end else if(T10) begin
      out_reg_9 <= io_in_11;
    end else if(T4) begin
      out_reg_9 <= io_in_9;
    end
    if(T14) begin
      out_reg_10 <= io_in_0;
    end else if(T12) begin
      out_reg_10 <= io_in_14;
    end else if(T10) begin
      out_reg_10 <= io_in_12;
    end else if(T4) begin
      out_reg_10 <= io_in_10;
    end
    if(T14) begin
      out_reg_11 <= io_in_1;
    end else if(T12) begin
      out_reg_11 <= io_in_15;
    end else if(T10) begin
      out_reg_11 <= io_in_13;
    end else if(T4) begin
      out_reg_11 <= io_in_11;
    end
    if(T14) begin
      out_reg_12 <= io_in_2;
    end else if(T12) begin
      out_reg_12 <= io_in_0;
    end else if(T10) begin
      out_reg_12 <= io_in_14;
    end else if(T4) begin
      out_reg_12 <= io_in_12;
    end
    if(T14) begin
      out_reg_13 <= io_in_3;
    end else if(T12) begin
      out_reg_13 <= io_in_1;
    end else if(T10) begin
      out_reg_13 <= io_in_15;
    end else if(T4) begin
      out_reg_13 <= io_in_13;
    end
    if(T14) begin
      out_reg_14 <= io_in_4;
    end else if(T12) begin
      out_reg_14 <= io_in_2;
    end else if(T10) begin
      out_reg_14 <= io_in_0;
    end else if(T4) begin
      out_reg_14 <= io_in_14;
    end
    if(T14) begin
      out_reg_15 <= io_in_5;
    end else if(T12) begin
      out_reg_15 <= io_in_3;
    end else if(T10) begin
      out_reg_15 <= io_in_1;
    end else if(T4) begin
      out_reg_15 <= io_in_15;
    end
    if(reset) begin
      start_next_stage_reg <= 1'h0;
    end else if(T8) begin
      start_next_stage_reg <= 1'h1;
    end
  end
endmodule

module streamMatrixTransposeTop(input clk, input reset,
    input  io_clk_en,
    input  io_start,
    output io_start_next_stage,
    input [63:0] io_in_15,
    input [63:0] io_in_14,
    input [63:0] io_in_13,
    input [63:0] io_in_12,
    input [63:0] io_in_11,
    input [63:0] io_in_10,
    input [63:0] io_in_9,
    input [63:0] io_in_8,
    input [63:0] io_in_7,
    input [63:0] io_in_6,
    input [63:0] io_in_5,
    input [63:0] io_in_4,
    input [63:0] io_in_3,
    input [63:0] io_in_2,
    input [63:0] io_in_1,
    input [63:0] io_in_0,
    output[63:0] io_out_15,
    output[63:0] io_out_14,
    output[63:0] io_out_13,
    output[63:0] io_out_12,
    output[63:0] io_out_11,
    output[63:0] io_out_10,
    output[63:0] io_out_9,
    output[63:0] io_out_8,
    output[63:0] io_out_7,
    output[63:0] io_out_6,
    output[63:0] io_out_5,
    output[63:0] io_out_4,
    output[63:0] io_out_3,
    output[63:0] io_out_2,
    output[63:0] io_out_1,
    output[63:0] io_out_0
);

  wire crossbar_io_start_next_stage;
  wire[63:0] crossbar_io_out_15;
  wire[63:0] crossbar_io_out_14;
  wire[63:0] crossbar_io_out_13;
  wire[63:0] crossbar_io_out_12;
  wire[63:0] crossbar_io_out_11;
  wire[63:0] crossbar_io_out_10;
  wire[63:0] crossbar_io_out_9;
  wire[63:0] crossbar_io_out_8;
  wire[63:0] crossbar_io_out_7;
  wire[63:0] crossbar_io_out_6;
  wire[63:0] crossbar_io_out_5;
  wire[63:0] crossbar_io_out_4;
  wire[63:0] crossbar_io_out_3;
  wire[63:0] crossbar_io_out_2;
  wire[63:0] crossbar_io_out_1;
  wire[63:0] crossbar_io_out_0;
  wire crossbarShift_io_start_next_stage;
  wire[63:0] crossbarShift_io_out_15;
  wire[63:0] crossbarShift_io_out_14;
  wire[63:0] crossbarShift_io_out_13;
  wire[63:0] crossbarShift_io_out_12;
  wire[63:0] crossbarShift_io_out_11;
  wire[63:0] crossbarShift_io_out_10;
  wire[63:0] crossbarShift_io_out_9;
  wire[63:0] crossbarShift_io_out_8;
  wire[63:0] crossbarShift_io_out_7;
  wire[63:0] crossbarShift_io_out_6;
  wire[63:0] crossbarShift_io_out_5;
  wire[63:0] crossbarShift_io_out_4;
  wire[63:0] crossbarShift_io_out_3;
  wire[63:0] crossbarShift_io_out_2;
  wire[63:0] crossbarShift_io_out_1;
  wire[63:0] crossbarShift_io_out_0;
  wire crossbarShift_1_io_start_next_stage;
  wire[63:0] crossbarShift_1_io_out_15;
  wire[63:0] crossbarShift_1_io_out_14;
  wire[63:0] crossbarShift_1_io_out_13;
  wire[63:0] crossbarShift_1_io_out_12;
  wire[63:0] crossbarShift_1_io_out_11;
  wire[63:0] crossbarShift_1_io_out_10;
  wire[63:0] crossbarShift_1_io_out_9;
  wire[63:0] crossbarShift_1_io_out_8;
  wire[63:0] crossbarShift_1_io_out_7;
  wire[63:0] crossbarShift_1_io_out_6;
  wire[63:0] crossbarShift_1_io_out_5;
  wire[63:0] crossbarShift_1_io_out_4;
  wire[63:0] crossbarShift_1_io_out_3;
  wire[63:0] crossbarShift_1_io_out_2;
  wire[63:0] crossbarShift_1_io_out_1;
  wire[63:0] crossbarShift_1_io_out_0;
  wire memArray_io_start_next_stage;
  wire[63:0] memArray_io_out_15;
  wire[63:0] memArray_io_out_14;
  wire[63:0] memArray_io_out_13;
  wire[63:0] memArray_io_out_12;
  wire[63:0] memArray_io_out_11;
  wire[63:0] memArray_io_out_10;
  wire[63:0] memArray_io_out_9;
  wire[63:0] memArray_io_out_8;
  wire[63:0] memArray_io_out_7;
  wire[63:0] memArray_io_out_6;
  wire[63:0] memArray_io_out_5;
  wire[63:0] memArray_io_out_4;
  wire[63:0] memArray_io_out_3;
  wire[63:0] memArray_io_out_2;
  wire[63:0] memArray_io_out_1;
  wire[63:0] memArray_io_out_0;


  assign io_out_0 = crossbarShift_1_io_out_0;
  assign io_out_1 = crossbarShift_1_io_out_1;
  assign io_out_2 = crossbarShift_1_io_out_2;
  assign io_out_3 = crossbarShift_1_io_out_3;
  assign io_out_4 = crossbarShift_1_io_out_4;
  assign io_out_5 = crossbarShift_1_io_out_5;
  assign io_out_6 = crossbarShift_1_io_out_6;
  assign io_out_7 = crossbarShift_1_io_out_7;
  assign io_out_8 = crossbarShift_1_io_out_8;
  assign io_out_9 = crossbarShift_1_io_out_9;
  assign io_out_10 = crossbarShift_1_io_out_10;
  assign io_out_11 = crossbarShift_1_io_out_11;
  assign io_out_12 = crossbarShift_1_io_out_12;
  assign io_out_13 = crossbarShift_1_io_out_13;
  assign io_out_14 = crossbarShift_1_io_out_14;
  assign io_out_15 = crossbarShift_1_io_out_15;
  assign io_start_next_stage = crossbarShift_1_io_start_next_stage;
  crossbar crossbar(.clk(clk), .reset(reset),
       .io_clk_en( io_clk_en ),
       .io_start( io_start ),
       .io_start_next_stage( crossbar_io_start_next_stage ),
       .io_in_15( io_in_15 ),
       .io_in_14( io_in_14 ),
       .io_in_13( io_in_13 ),
       .io_in_12( io_in_12 ),
       .io_in_11( io_in_11 ),
       .io_in_10( io_in_10 ),
       .io_in_9( io_in_9 ),
       .io_in_8( io_in_8 ),
       .io_in_7( io_in_7 ),
       .io_in_6( io_in_6 ),
       .io_in_5( io_in_5 ),
       .io_in_4( io_in_4 ),
       .io_in_3( io_in_3 ),
       .io_in_2( io_in_2 ),
       .io_in_1( io_in_1 ),
       .io_in_0( io_in_0 ),
       .io_out_15( crossbar_io_out_15 ),
       .io_out_14( crossbar_io_out_14 ),
       .io_out_13( crossbar_io_out_13 ),
       .io_out_12( crossbar_io_out_12 ),
       .io_out_11( crossbar_io_out_11 ),
       .io_out_10( crossbar_io_out_10 ),
       .io_out_9( crossbar_io_out_9 ),
       .io_out_8( crossbar_io_out_8 ),
       .io_out_7( crossbar_io_out_7 ),
       .io_out_6( crossbar_io_out_6 ),
       .io_out_5( crossbar_io_out_5 ),
       .io_out_4( crossbar_io_out_4 ),
       .io_out_3( crossbar_io_out_3 ),
       .io_out_2( crossbar_io_out_2 ),
       .io_out_1( crossbar_io_out_1 ),
       .io_out_0( crossbar_io_out_0 )
  );
  crossbarShiftDown crossbarShift(.clk(clk), .reset(reset),
       .io_clk_en( io_clk_en ),
       .io_start( crossbar_io_start_next_stage ),
       .io_start_next_stage( crossbarShift_io_start_next_stage ),
       .io_in_15( crossbar_io_out_15 ),
       .io_in_14( crossbar_io_out_14 ),
       .io_in_13( crossbar_io_out_13 ),
       .io_in_12( crossbar_io_out_12 ),
       .io_in_11( crossbar_io_out_11 ),
       .io_in_10( crossbar_io_out_10 ),
       .io_in_9( crossbar_io_out_9 ),
       .io_in_8( crossbar_io_out_8 ),
       .io_in_7( crossbar_io_out_7 ),
       .io_in_6( crossbar_io_out_6 ),
       .io_in_5( crossbar_io_out_5 ),
       .io_in_4( crossbar_io_out_4 ),
       .io_in_3( crossbar_io_out_3 ),
       .io_in_2( crossbar_io_out_2 ),
       .io_in_1( crossbar_io_out_1 ),
       .io_in_0( crossbar_io_out_0 ),
       .io_out_15( crossbarShift_io_out_15 ),
       .io_out_14( crossbarShift_io_out_14 ),
       .io_out_13( crossbarShift_io_out_13 ),
       .io_out_12( crossbarShift_io_out_12 ),
       .io_out_11( crossbarShift_io_out_11 ),
       .io_out_10( crossbarShift_io_out_10 ),
       .io_out_9( crossbarShift_io_out_9 ),
       .io_out_8( crossbarShift_io_out_8 ),
       .io_out_7( crossbarShift_io_out_7 ),
       .io_out_6( crossbarShift_io_out_6 ),
       .io_out_5( crossbarShift_io_out_5 ),
       .io_out_4( crossbarShift_io_out_4 ),
       .io_out_3( crossbarShift_io_out_3 ),
       .io_out_2( crossbarShift_io_out_2 ),
       .io_out_1( crossbarShift_io_out_1 ),
       .io_out_0( crossbarShift_io_out_0 )
  );
  memArray memArray(.clk(clk), .reset(reset),
       .io_clk_en( io_clk_en ),
       .io_start( crossbarShift_io_start_next_stage ),
       .io_start_next_stage( memArray_io_start_next_stage ),
       .io_in_15( crossbarShift_io_out_15 ),
       .io_in_14( crossbarShift_io_out_14 ),
       .io_in_13( crossbarShift_io_out_13 ),
       .io_in_12( crossbarShift_io_out_12 ),
       .io_in_11( crossbarShift_io_out_11 ),
       .io_in_10( crossbarShift_io_out_10 ),
       .io_in_9( crossbarShift_io_out_9 ),
       .io_in_8( crossbarShift_io_out_8 ),
       .io_in_7( crossbarShift_io_out_7 ),
       .io_in_6( crossbarShift_io_out_6 ),
       .io_in_5( crossbarShift_io_out_5 ),
       .io_in_4( crossbarShift_io_out_4 ),
       .io_in_3( crossbarShift_io_out_3 ),
       .io_in_2( crossbarShift_io_out_2 ),
       .io_in_1( crossbarShift_io_out_1 ),
       .io_in_0( crossbarShift_io_out_0 ),
       .io_out_15( memArray_io_out_15 ),
       .io_out_14( memArray_io_out_14 ),
       .io_out_13( memArray_io_out_13 ),
       .io_out_12( memArray_io_out_12 ),
       .io_out_11( memArray_io_out_11 ),
       .io_out_10( memArray_io_out_10 ),
       .io_out_9( memArray_io_out_9 ),
       .io_out_8( memArray_io_out_8 ),
       .io_out_7( memArray_io_out_7 ),
       .io_out_6( memArray_io_out_6 ),
       .io_out_5( memArray_io_out_5 ),
       .io_out_4( memArray_io_out_4 ),
       .io_out_3( memArray_io_out_3 ),
       .io_out_2( memArray_io_out_2 ),
       .io_out_1( memArray_io_out_1 ),
       .io_out_0( memArray_io_out_0 )
  );
  crossbarShiftUp crossbarShift_1(.clk(clk), .reset(reset),
       .io_clk_en( io_clk_en ),
       .io_start( memArray_io_start_next_stage ),
       .io_start_next_stage( crossbarShift_1_io_start_next_stage ),
       .io_in_15( memArray_io_out_15 ),
       .io_in_14( memArray_io_out_14 ),
       .io_in_13( memArray_io_out_13 ),
       .io_in_12( memArray_io_out_12 ),
       .io_in_11( memArray_io_out_11 ),
       .io_in_10( memArray_io_out_10 ),
       .io_in_9( memArray_io_out_9 ),
       .io_in_8( memArray_io_out_8 ),
       .io_in_7( memArray_io_out_7 ),
       .io_in_6( memArray_io_out_6 ),
       .io_in_5( memArray_io_out_5 ),
       .io_in_4( memArray_io_out_4 ),
       .io_in_3( memArray_io_out_3 ),
       .io_in_2( memArray_io_out_2 ),
       .io_in_1( memArray_io_out_1 ),
       .io_in_0( memArray_io_out_0 ),
       .io_out_15( crossbarShift_1_io_out_15 ),
       .io_out_14( crossbarShift_1_io_out_14 ),
       .io_out_13( crossbarShift_1_io_out_13 ),
       .io_out_12( crossbarShift_1_io_out_12 ),
       .io_out_11( crossbarShift_1_io_out_11 ),
       .io_out_10( crossbarShift_1_io_out_10 ),
       .io_out_9( crossbarShift_1_io_out_9 ),
       .io_out_8( crossbarShift_1_io_out_8 ),
       .io_out_7( crossbarShift_1_io_out_7 ),
       .io_out_6( crossbarShift_1_io_out_6 ),
       .io_out_5( crossbarShift_1_io_out_5 ),
       .io_out_4( crossbarShift_1_io_out_4 ),
       .io_out_3( crossbarShift_1_io_out_3 ),
       .io_out_2( crossbarShift_1_io_out_2 ),
       .io_out_1( crossbarShift_1_io_out_1 ),
       .io_out_0( crossbarShift_1_io_out_0 )
  );
endmodule

module multComplex(input clk, input reset,
    input [31:0] io_real1,
    input [31:0] io_img1,
    input [31:0] io_real2,
    input [31:0] io_img2,
    output[31:0] io_realOut,
    output[31:0] io_imgOut
);

  reg [31:0] delayArrayReal1_1;
  reg [31:0] delayArrayReal1_0;
  reg [31:0] delayArrayImg1_1;
  reg [31:0] delayArrayImg1_0;
  reg [31:0] delayArrayReal2_1;
  reg [31:0] delayArrayReal2_0;
  wire[31:0] addsubfxp_q;
  wire[31:0] addsubfxp_1_q;
  wire[31:0] addsubfxp_2_q;
  wire[31:0] addsubfxp_3_q;
  wire[31:0] addsubfxp_4_q;
  wire[31:0] multfix_q_sc;
  wire[31:0] multfix_1_q_sc;
  wire[31:0] multfix_2_q_sc;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    delayArrayReal1_1 = {1{$random}};
    delayArrayReal1_0 = {1{$random}};
    delayArrayImg1_1 = {1{$random}};
    delayArrayImg1_0 = {1{$random}};
    delayArrayReal2_1 = {1{$random}};
    delayArrayReal2_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_imgOut = addsubfxp_2_q;
  assign io_realOut = addsubfxp_4_q;
  subfxp # (
    .width(32),
    .cycles(2)
  ) addsubfxp(.clk(clk),
       .a( io_real1 ),
       .b( io_img1 ),
       .q( addsubfxp_q )
  );
  subfxp # (
    .width(32),
    .cycles(2)
  ) addsubfxp_1(.clk(clk),
       .a( io_real2 ),
       .b( io_img2 ),
       .q( addsubfxp_1_q )
  );
  subfxp # (
    .width(32),
    .cycles(2)
  ) addsubfxp_2(.clk(clk),
       .a( multfix_q_sc ),
       .b( multfix_2_q_sc ),
       .q( addsubfxp_2_q )
  );
  addfxp # (
    .width(32),
    .cycles(2)
  ) addsubfxp_3(.clk(clk),
       .a( io_real2 ),
       .b( io_img2 ),
       .q( addsubfxp_3_q )
  );
  addfxp # (
    .width(32),
    .cycles(2)
  ) addsubfxp_4(.clk(clk),
       .a( multfix_q_sc ),
       .b( multfix_1_q_sc ),
       .q( addsubfxp_4_q )
  );
  multfix # (
    .WIDTH(32),
    .CYCLES(1)
  ) multfix(.clk(clk), .rst(reset),
       .a( addsubfxp_q ),
       .b( delayArrayReal2_1 ),
       .q_sc( multfix_q_sc )
       //.q_unsc(  )
  );
  multfix # (
    .WIDTH(32),
    .CYCLES(1)
  ) multfix_1(.clk(clk), .rst(reset),
       .a( delayArrayImg1_1 ),
       .b( addsubfxp_1_q ),
       .q_sc( multfix_1_q_sc )
       //.q_unsc(  )
  );
  multfix # (
    .WIDTH(32),
    .CYCLES(1)
  ) multfix_2(.clk(clk), .rst(reset),
       .a( addsubfxp_3_q ),
       .b( delayArrayReal1_1 ),
       .q_sc( multfix_2_q_sc )
       //.q_unsc(  )
  );

  always @(posedge clk) begin
    delayArrayReal1_1 <= delayArrayReal1_0;
    delayArrayReal1_0 <= io_real1;
    delayArrayImg1_1 <= delayArrayImg1_0;
    delayArrayImg1_0 <= io_img1;
    delayArrayReal2_1 <= delayArrayReal2_0;
    delayArrayReal2_0 <= io_real2;
  end
endmodule

module two_d_convolution(input clk, input reset,
    input  io_clk_en,
    input  io_start,
    output io_start_next_stage,
    input [31:0] io_in_15,
    input [31:0] io_in_14,
    input [31:0] io_in_13,
    input [31:0] io_in_12,
    input [31:0] io_in_11,
    input [31:0] io_in_10,
    input [31:0] io_in_9,
    input [31:0] io_in_8,
    input [31:0] io_in_7,
    input [31:0] io_in_6,
    input [31:0] io_in_5,
    input [31:0] io_in_4,
    input [31:0] io_in_3,
    input [31:0] io_in_2,
    input [31:0] io_in_1,
    input [31:0] io_in_0,
    output[31:0] io_out_15,
    output[31:0] io_out_14,
    output[31:0] io_out_13,
    output[31:0] io_out_12,
    output[31:0] io_out_11,
    output[31:0] io_out_10,
    output[31:0] io_out_9,
    output[31:0] io_out_8,
    output[31:0] io_out_7,
    output[31:0] io_out_6,
    output[31:0] io_out_5,
    output[31:0] io_out_4,
    output[31:0] io_out_3,
    output[31:0] io_out_2,
    output[31:0] io_out_1,
    output[31:0] io_out_0
);

  wire[63:0] T0;
  wire[63:0] T1;
  wire[63:0] T2;
  wire[63:0] T3;
  wire[63:0] T4;
  wire[63:0] T5;
  wire[63:0] T6;
  wire[63:0] T7;
  wire[63:0] T8;
  wire[63:0] T9;
  wire[63:0] T10;
  wire[63:0] T11;
  wire[63:0] T12;
  wire[63:0] T13;
  wire[63:0] T14;
  wire[63:0] T15;
  reg  startSecondMatrix;
  wire[31:0] T16;
  reg [63:0] delaySecond_8;
  wire[31:0] T17;
  wire[31:0] T18;
  reg [63:0] delaySecond_9;
  wire[31:0] T19;
  wire[31:0] T20;
  reg [63:0] delaySecond_10;
  wire[31:0] T21;
  wire[31:0] T22;
  reg [63:0] delaySecond_11;
  wire[31:0] T23;
  wire[31:0] T24;
  reg [63:0] delaySecond_12;
  wire[31:0] T25;
  wire[31:0] T26;
  reg [63:0] delaySecond_13;
  wire[31:0] T27;
  wire[31:0] T28;
  reg [63:0] delaySecond_14;
  wire[31:0] T29;
  wire[31:0] T30;
  reg [63:0] delaySecond_15;
  wire[31:0] T31;
  wire[31:0] T32;
  reg [63:0] delaySecond_0;
  wire[31:0] T33;
  wire[31:0] T34;
  reg [63:0] delaySecond_1;
  wire[31:0] T35;
  wire[31:0] T36;
  reg [63:0] delaySecond_2;
  wire[31:0] T37;
  wire[31:0] T38;
  reg [63:0] delaySecond_3;
  wire[31:0] T39;
  wire[31:0] T40;
  reg [63:0] delaySecond_4;
  wire[31:0] T41;
  wire[31:0] T42;
  reg [63:0] delaySecond_5;
  wire[31:0] T43;
  wire[31:0] T44;
  reg [63:0] delaySecond_6;
  wire[31:0] T45;
  wire[31:0] T46;
  reg [63:0] delaySecond_7;
  wire[31:0] T47;
  reg  delayArrayNext_2;
  reg  delayArrayNext_1;
  reg  delayArrayNext_0;
  wire[31:0] T48;
  reg [63:0] delayFirst_8;
  wire[31:0] T49;
  wire[31:0] T50;
  reg [63:0] delayFirst_9;
  wire[31:0] T51;
  wire[31:0] T52;
  reg [63:0] delayFirst_10;
  wire[31:0] T53;
  wire[31:0] T54;
  reg [63:0] delayFirst_11;
  wire[31:0] T55;
  wire[31:0] T56;
  reg [63:0] delayFirst_12;
  wire[31:0] T57;
  wire[31:0] T58;
  reg [63:0] delayFirst_13;
  wire[31:0] T59;
  wire[31:0] T60;
  reg [63:0] delayFirst_14;
  wire[31:0] T61;
  wire[31:0] T62;
  reg [63:0] delayFirst_15;
  wire[31:0] T63;
  wire[31:0] T64;
  reg [63:0] delayFirst_0;
  wire[31:0] T65;
  wire[31:0] T66;
  reg [63:0] delayFirst_1;
  wire[31:0] T67;
  wire[31:0] T68;
  reg [63:0] delayFirst_2;
  wire[31:0] T69;
  wire[31:0] T70;
  reg [63:0] delayFirst_3;
  wire[31:0] T71;
  wire[31:0] T72;
  reg [63:0] delayFirst_4;
  wire[31:0] T73;
  wire[31:0] T74;
  reg [63:0] delayFirst_5;
  wire[31:0] T75;
  wire[31:0] T76;
  reg [63:0] delayFirst_6;
  wire[31:0] T77;
  wire[31:0] T78;
  reg [63:0] delayFirst_7;
  wire[31:0] T79;
  wire[63:0] T80;
  wire[63:0] T81;
  wire[63:0] T82;
  wire[63:0] T83;
  wire[63:0] T84;
  wire[63:0] T85;
  wire[63:0] T86;
  wire[63:0] T87;
  wire[63:0] T88;
  wire[63:0] T89;
  wire[63:0] T90;
  wire[63:0] T91;
  wire[63:0] T92;
  wire[63:0] T93;
  wire[63:0] T94;
  wire[63:0] T95;
  reg  startFirstMatrix;
  reg [31:0] delayInput_8;
  reg [31:0] delayInput_9;
  reg [31:0] delayInput_10;
  reg [31:0] delayInput_11;
  reg [31:0] delayInput_12;
  reg [31:0] delayInput_13;
  reg [31:0] delayInput_14;
  reg [31:0] delayInput_15;
  reg [31:0] delayInput_0;
  reg [31:0] delayInput_1;
  reg [31:0] delayInput_2;
  reg [31:0] delayInput_3;
  reg [31:0] delayInput_4;
  reg [31:0] delayInput_5;
  reg [31:0] delayInput_6;
  reg [31:0] delayInput_7;
  reg  delayStartNextStage;
  wire fft_next_out;
  wire[31:0] fft_Y15;
  wire[31:0] fft_Y14;
  wire[31:0] fft_Y13;
  wire[31:0] fft_Y12;
  wire[31:0] fft_Y11;
  wire[31:0] fft_Y10;
  wire[31:0] fft_Y9;
  wire[31:0] fft_Y8;
  wire[31:0] fft_Y7;
  wire[31:0] fft_Y6;
  wire[31:0] fft_Y5;
  wire[31:0] fft_Y4;
  wire[31:0] fft_Y3;
  wire[31:0] fft_Y2;
  wire[31:0] fft_Y1;
  wire[31:0] fft_Y0;
  wire[31:0] fft_1_Y15;
  wire[31:0] fft_1_Y14;
  wire[31:0] fft_1_Y13;
  wire[31:0] fft_1_Y12;
  wire[31:0] fft_1_Y11;
  wire[31:0] fft_1_Y10;
  wire[31:0] fft_1_Y9;
  wire[31:0] fft_1_Y8;
  wire[31:0] fft_1_Y7;
  wire[31:0] fft_1_Y6;
  wire[31:0] fft_1_Y5;
  wire[31:0] fft_1_Y4;
  wire[31:0] fft_1_Y3;
  wire[31:0] fft_1_Y2;
  wire[31:0] fft_1_Y1;
  wire[31:0] fft_1_Y0;
  wire fft_2_next_out;
  wire[31:0] fft_2_Y15;
  wire[31:0] fft_2_Y14;
  wire[31:0] fft_2_Y13;
  wire[31:0] fft_2_Y12;
  wire[31:0] fft_2_Y11;
  wire[31:0] fft_2_Y10;
  wire[31:0] fft_2_Y9;
  wire[31:0] fft_2_Y8;
  wire[31:0] fft_2_Y7;
  wire[31:0] fft_2_Y6;
  wire[31:0] fft_2_Y5;
  wire[31:0] fft_2_Y4;
  wire[31:0] fft_2_Y3;
  wire[31:0] fft_2_Y2;
  wire[31:0] fft_2_Y1;
  wire[31:0] fft_2_Y0;
  wire[31:0] fft_3_Y15;
  wire[31:0] fft_3_Y14;
  wire[31:0] fft_3_Y13;
  wire[31:0] fft_3_Y12;
  wire[31:0] fft_3_Y11;
  wire[31:0] fft_3_Y10;
  wire[31:0] fft_3_Y9;
  wire[31:0] fft_3_Y8;
  wire[31:0] fft_3_Y7;
  wire[31:0] fft_3_Y6;
  wire[31:0] fft_3_Y5;
  wire[31:0] fft_3_Y4;
  wire[31:0] fft_3_Y3;
  wire[31:0] fft_3_Y2;
  wire[31:0] fft_3_Y1;
  wire[31:0] fft_3_Y0;
  wire fft_4_next_out;
  wire[31:0] fft_4_Y15;
  wire[31:0] fft_4_Y14;
  wire[31:0] fft_4_Y13;
  wire[31:0] fft_4_Y12;
  wire[31:0] fft_4_Y11;
  wire[31:0] fft_4_Y10;
  wire[31:0] fft_4_Y9;
  wire[31:0] fft_4_Y8;
  wire[31:0] fft_4_Y7;
  wire[31:0] fft_4_Y6;
  wire[31:0] fft_4_Y5;
  wire[31:0] fft_4_Y4;
  wire[31:0] fft_4_Y3;
  wire[31:0] fft_4_Y2;
  wire[31:0] fft_4_Y1;
  wire[31:0] fft_4_Y0;
  wire[31:0] fft_5_Y15;
  wire[31:0] fft_5_Y14;
  wire[31:0] fft_5_Y13;
  wire[31:0] fft_5_Y12;
  wire[31:0] fft_5_Y11;
  wire[31:0] fft_5_Y10;
  wire[31:0] fft_5_Y9;
  wire[31:0] fft_5_Y8;
  wire[31:0] fft_5_Y7;
  wire[31:0] fft_5_Y6;
  wire[31:0] fft_5_Y5;
  wire[31:0] fft_5_Y4;
  wire[31:0] fft_5_Y3;
  wire[31:0] fft_5_Y2;
  wire[31:0] fft_5_Y1;
  wire[31:0] fft_5_Y0;
  wire fft_6_next_out;
  wire[31:0] fft_6_Y14;
  wire[31:0] fft_6_Y12;
  wire[31:0] fft_6_Y10;
  wire[31:0] fft_6_Y8;
  wire[31:0] fft_6_Y6;
  wire[31:0] fft_6_Y4;
  wire[31:0] fft_6_Y2;
  wire[31:0] fft_6_Y0;
  wire[31:0] fft_7_Y14;
  wire[31:0] fft_7_Y12;
  wire[31:0] fft_7_Y10;
  wire[31:0] fft_7_Y8;
  wire[31:0] fft_7_Y6;
  wire[31:0] fft_7_Y4;
  wire[31:0] fft_7_Y2;
  wire[31:0] fft_7_Y0;
  wire[31:0] multComplex_io_realOut;
  wire[31:0] multComplex_io_imgOut;
  wire[31:0] multComplex_1_io_realOut;
  wire[31:0] multComplex_1_io_imgOut;
  wire[31:0] multComplex_2_io_realOut;
  wire[31:0] multComplex_2_io_imgOut;
  wire[31:0] multComplex_3_io_realOut;
  wire[31:0] multComplex_3_io_imgOut;
  wire[31:0] multComplex_4_io_realOut;
  wire[31:0] multComplex_4_io_imgOut;
  wire[31:0] multComplex_5_io_realOut;
  wire[31:0] multComplex_5_io_imgOut;
  wire[31:0] multComplex_6_io_realOut;
  wire[31:0] multComplex_6_io_imgOut;
  wire[31:0] multComplex_7_io_realOut;
  wire[31:0] multComplex_7_io_imgOut;
  wire[31:0] multComplex_8_io_realOut;
  wire[31:0] multComplex_8_io_imgOut;
  wire[31:0] multComplex_9_io_realOut;
  wire[31:0] multComplex_9_io_imgOut;
  wire[31:0] multComplex_10_io_realOut;
  wire[31:0] multComplex_10_io_imgOut;
  wire[31:0] multComplex_11_io_realOut;
  wire[31:0] multComplex_11_io_imgOut;
  wire[31:0] multComplex_12_io_realOut;
  wire[31:0] multComplex_12_io_imgOut;
  wire[31:0] multComplex_13_io_realOut;
  wire[31:0] multComplex_13_io_imgOut;
  wire[31:0] multComplex_14_io_realOut;
  wire[31:0] multComplex_14_io_imgOut;
  wire[31:0] multComplex_15_io_realOut;
  wire[31:0] multComplex_15_io_imgOut;
  wire streamMatrixTransposeTop_io_start_next_stage;
  wire[63:0] streamMatrixTransposeTop_io_out_15;
  wire[63:0] streamMatrixTransposeTop_io_out_14;
  wire[63:0] streamMatrixTransposeTop_io_out_13;
  wire[63:0] streamMatrixTransposeTop_io_out_12;
  wire[63:0] streamMatrixTransposeTop_io_out_11;
  wire[63:0] streamMatrixTransposeTop_io_out_10;
  wire[63:0] streamMatrixTransposeTop_io_out_9;
  wire[63:0] streamMatrixTransposeTop_io_out_8;
  wire[63:0] streamMatrixTransposeTop_io_out_7;
  wire[63:0] streamMatrixTransposeTop_io_out_6;
  wire[63:0] streamMatrixTransposeTop_io_out_5;
  wire[63:0] streamMatrixTransposeTop_io_out_4;
  wire[63:0] streamMatrixTransposeTop_io_out_3;
  wire[63:0] streamMatrixTransposeTop_io_out_2;
  wire[63:0] streamMatrixTransposeTop_io_out_1;
  wire[63:0] streamMatrixTransposeTop_io_out_0;
  wire streamMatrixTransposeTop_1_io_start_next_stage;
  wire[63:0] streamMatrixTransposeTop_1_io_out_15;
  wire[63:0] streamMatrixTransposeTop_1_io_out_14;
  wire[63:0] streamMatrixTransposeTop_1_io_out_13;
  wire[63:0] streamMatrixTransposeTop_1_io_out_12;
  wire[63:0] streamMatrixTransposeTop_1_io_out_11;
  wire[63:0] streamMatrixTransposeTop_1_io_out_10;
  wire[63:0] streamMatrixTransposeTop_1_io_out_9;
  wire[63:0] streamMatrixTransposeTop_1_io_out_8;
  wire[63:0] streamMatrixTransposeTop_1_io_out_7;
  wire[63:0] streamMatrixTransposeTop_1_io_out_6;
  wire[63:0] streamMatrixTransposeTop_1_io_out_5;
  wire[63:0] streamMatrixTransposeTop_1_io_out_4;
  wire[63:0] streamMatrixTransposeTop_1_io_out_3;
  wire[63:0] streamMatrixTransposeTop_1_io_out_2;
  wire[63:0] streamMatrixTransposeTop_1_io_out_1;
  wire[63:0] streamMatrixTransposeTop_1_io_out_0;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    startSecondMatrix = {1{$random}};
    delaySecond_8 = {2{$random}};
    delaySecond_9 = {2{$random}};
    delaySecond_10 = {2{$random}};
    delaySecond_11 = {2{$random}};
    delaySecond_12 = {2{$random}};
    delaySecond_13 = {2{$random}};
    delaySecond_14 = {2{$random}};
    delaySecond_15 = {2{$random}};
    delaySecond_0 = {2{$random}};
    delaySecond_1 = {2{$random}};
    delaySecond_2 = {2{$random}};
    delaySecond_3 = {2{$random}};
    delaySecond_4 = {2{$random}};
    delaySecond_5 = {2{$random}};
    delaySecond_6 = {2{$random}};
    delaySecond_7 = {2{$random}};
    delayArrayNext_2 = {1{$random}};
    delayArrayNext_1 = {1{$random}};
    delayArrayNext_0 = {1{$random}};
    delayFirst_8 = {2{$random}};
    delayFirst_9 = {2{$random}};
    delayFirst_10 = {2{$random}};
    delayFirst_11 = {2{$random}};
    delayFirst_12 = {2{$random}};
    delayFirst_13 = {2{$random}};
    delayFirst_14 = {2{$random}};
    delayFirst_15 = {2{$random}};
    delayFirst_0 = {2{$random}};
    delayFirst_1 = {2{$random}};
    delayFirst_2 = {2{$random}};
    delayFirst_3 = {2{$random}};
    delayFirst_4 = {2{$random}};
    delayFirst_5 = {2{$random}};
    delayFirst_6 = {2{$random}};
    delayFirst_7 = {2{$random}};
    startFirstMatrix = {1{$random}};
    delayInput_8 = {1{$random}};
    delayInput_9 = {1{$random}};
    delayInput_10 = {1{$random}};
    delayInput_11 = {1{$random}};
    delayInput_12 = {1{$random}};
    delayInput_13 = {1{$random}};
    delayInput_14 = {1{$random}};
    delayInput_15 = {1{$random}};
    delayInput_0 = {1{$random}};
    delayInput_1 = {1{$random}};
    delayInput_2 = {1{$random}};
    delayInput_3 = {1{$random}};
    delayInput_4 = {1{$random}};
    delayInput_5 = {1{$random}};
    delayInput_6 = {1{$random}};
    delayInput_7 = {1{$random}};
    delayStartNextStage = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = {fft_4_Y1, fft_4_Y0};
  assign T1 = {fft_4_Y3, fft_4_Y2};
  assign T2 = {fft_4_Y5, fft_4_Y4};
  assign T3 = {fft_4_Y7, fft_4_Y6};
  assign T4 = {fft_4_Y9, fft_4_Y8};
  assign T5 = {fft_4_Y11, fft_4_Y10};
  assign T6 = {fft_4_Y13, fft_4_Y12};
  assign T7 = {fft_4_Y15, fft_4_Y14};
  assign T8 = {fft_5_Y1, fft_5_Y0};
  assign T9 = {fft_5_Y3, fft_5_Y2};
  assign T10 = {fft_5_Y5, fft_5_Y4};
  assign T11 = {fft_5_Y7, fft_5_Y6};
  assign T12 = {fft_5_Y9, fft_5_Y8};
  assign T13 = {fft_5_Y11, fft_5_Y10};
  assign T14 = {fft_5_Y13, fft_5_Y12};
  assign T15 = {fft_5_Y15, fft_5_Y14};
  assign T16 = delaySecond_8[31:0];
  assign T17 = delaySecond_8[63:32];
  assign T18 = delaySecond_9[31:0];
  assign T19 = delaySecond_9[63:32];
  assign T20 = delaySecond_10[31:0];
  assign T21 = delaySecond_10[63:32];
  assign T22 = delaySecond_11[31:0];
  assign T23 = delaySecond_11[63:32];
  assign T24 = delaySecond_12[31:0];
  assign T25 = delaySecond_12[63:32];
  assign T26 = delaySecond_13[31:0];
  assign T27 = delaySecond_13[63:32];
  assign T28 = delaySecond_14[31:0];
  assign T29 = delaySecond_14[63:32];
  assign T30 = delaySecond_15[31:0];
  assign T31 = delaySecond_15[63:32];
  assign T32 = delaySecond_0[31:0];
  assign T33 = delaySecond_0[63:32];
  assign T34 = delaySecond_1[31:0];
  assign T35 = delaySecond_1[63:32];
  assign T36 = delaySecond_2[31:0];
  assign T37 = delaySecond_2[63:32];
  assign T38 = delaySecond_3[31:0];
  assign T39 = delaySecond_3[63:32];
  assign T40 = delaySecond_4[31:0];
  assign T41 = delaySecond_4[63:32];
  assign T42 = delaySecond_5[31:0];
  assign T43 = delaySecond_5[63:32];
  assign T44 = delaySecond_6[31:0];
  assign T45 = delaySecond_6[63:32];
  assign T46 = delaySecond_7[31:0];
  assign T47 = delaySecond_7[63:32];
  assign T48 = delayFirst_8[31:0];
  assign T49 = delayFirst_8[63:32];
  assign T50 = delayFirst_9[31:0];
  assign T51 = delayFirst_9[63:32];
  assign T52 = delayFirst_10[31:0];
  assign T53 = delayFirst_10[63:32];
  assign T54 = delayFirst_11[31:0];
  assign T55 = delayFirst_11[63:32];
  assign T56 = delayFirst_12[31:0];
  assign T57 = delayFirst_12[63:32];
  assign T58 = delayFirst_13[31:0];
  assign T59 = delayFirst_13[63:32];
  assign T60 = delayFirst_14[31:0];
  assign T61 = delayFirst_14[63:32];
  assign T62 = delayFirst_15[31:0];
  assign T63 = delayFirst_15[63:32];
  assign T64 = delayFirst_0[31:0];
  assign T65 = delayFirst_0[63:32];
  assign T66 = delayFirst_1[31:0];
  assign T67 = delayFirst_1[63:32];
  assign T68 = delayFirst_2[31:0];
  assign T69 = delayFirst_2[63:32];
  assign T70 = delayFirst_3[31:0];
  assign T71 = delayFirst_3[63:32];
  assign T72 = delayFirst_4[31:0];
  assign T73 = delayFirst_4[63:32];
  assign T74 = delayFirst_5[31:0];
  assign T75 = delayFirst_5[63:32];
  assign T76 = delayFirst_6[31:0];
  assign T77 = delayFirst_6[63:32];
  assign T78 = delayFirst_7[31:0];
  assign T79 = delayFirst_7[63:32];
  assign T80 = {fft_Y1, fft_Y0};
  assign T81 = {fft_Y3, fft_Y2};
  assign T82 = {fft_Y5, fft_Y4};
  assign T83 = {fft_Y7, fft_Y6};
  assign T84 = {fft_Y9, fft_Y8};
  assign T85 = {fft_Y11, fft_Y10};
  assign T86 = {fft_Y13, fft_Y12};
  assign T87 = {fft_Y15, fft_Y14};
  assign T88 = {fft_1_Y1, fft_1_Y0};
  assign T89 = {fft_1_Y3, fft_1_Y2};
  assign T90 = {fft_1_Y5, fft_1_Y4};
  assign T91 = {fft_1_Y7, fft_1_Y6};
  assign T92 = {fft_1_Y9, fft_1_Y8};
  assign T93 = {fft_1_Y11, fft_1_Y10};
  assign T94 = {fft_1_Y13, fft_1_Y12};
  assign T95 = {fft_1_Y15, fft_1_Y14};
  assign io_out_0 = fft_6_Y0;
  assign io_out_1 = fft_6_Y2;
  assign io_out_2 = fft_6_Y4;
  assign io_out_3 = fft_6_Y6;
  assign io_out_4 = fft_6_Y8;
  assign io_out_5 = fft_6_Y10;
  assign io_out_6 = fft_6_Y12;
  assign io_out_7 = fft_6_Y14;
  assign io_out_8 = fft_7_Y0;
  assign io_out_9 = fft_7_Y2;
  assign io_out_10 = fft_7_Y4;
  assign io_out_11 = fft_7_Y6;
  assign io_out_12 = fft_7_Y8;
  assign io_out_13 = fft_7_Y10;
  assign io_out_14 = fft_7_Y12;
  assign io_out_15 = fft_7_Y14;
  assign io_start_next_stage = delayStartNextStage;
  fft8_8 fft(.clk(clk), .reset(reset),
       .next( io_start ),
       .next_out( fft_next_out ),
       .X15( 32'h0 ),
       .X14( delayInput_7 ),
       .X13( 32'h0 ),
       .X12( delayInput_6 ),
       .X11( 32'h0 ),
       .X10( delayInput_5 ),
       .X9( 32'h0 ),
       .X8( delayInput_4 ),
       .X7( 32'h0 ),
       .X6( delayInput_3 ),
       .X5( 32'h0 ),
       .X4( delayInput_2 ),
       .X3( 32'h0 ),
       .X2( delayInput_1 ),
       .X1( 32'h0 ),
       .X0( delayInput_0 ),
       .Y15( fft_Y15 ),
       .Y14( fft_Y14 ),
       .Y13( fft_Y13 ),
       .Y12( fft_Y12 ),
       .Y11( fft_Y11 ),
       .Y10( fft_Y10 ),
       .Y9( fft_Y9 ),
       .Y8( fft_Y8 ),
       .Y7( fft_Y7 ),
       .Y6( fft_Y6 ),
       .Y5( fft_Y5 ),
       .Y4( fft_Y4 ),
       .Y3( fft_Y3 ),
       .Y2( fft_Y2 ),
       .Y1( fft_Y1 ),
       .Y0( fft_Y0 )
  );
  fft8_8 fft_1(.clk(clk), .reset(reset),
       .next( io_start ),
       //.next_out(  )
       .X15( 32'h0 ),
       .X14( delayInput_15 ),
       .X13( 32'h0 ),
       .X12( delayInput_14 ),
       .X11( 32'h0 ),
       .X10( delayInput_13 ),
       .X9( 32'h0 ),
       .X8( delayInput_12 ),
       .X7( 32'h0 ),
       .X6( delayInput_11 ),
       .X5( 32'h0 ),
       .X4( delayInput_10 ),
       .X3( 32'h0 ),
       .X2( delayInput_9 ),
       .X1( 32'h0 ),
       .X0( delayInput_8 ),
       .Y15( fft_1_Y15 ),
       .Y14( fft_1_Y14 ),
       .Y13( fft_1_Y13 ),
       .Y12( fft_1_Y12 ),
       .Y11( fft_1_Y11 ),
       .Y10( fft_1_Y10 ),
       .Y9( fft_1_Y9 ),
       .Y8( fft_1_Y8 ),
       .Y7( fft_1_Y7 ),
       .Y6( fft_1_Y6 ),
       .Y5( fft_1_Y5 ),
       .Y4( fft_1_Y4 ),
       .Y3( fft_1_Y3 ),
       .Y2( fft_1_Y2 ),
       .Y1( fft_1_Y1 ),
       .Y0( fft_1_Y0 )
  );
  streamMatrixTransposeTop streamMatrixTransposeTop(.clk(clk), .reset(reset),
       .io_clk_en( 1'h1 ),
       .io_start( startFirstMatrix ),
       .io_start_next_stage( streamMatrixTransposeTop_io_start_next_stage ),
       .io_in_15( T95 ),
       .io_in_14( T94 ),
       .io_in_13( T93 ),
       .io_in_12( T92 ),
       .io_in_11( T91 ),
       .io_in_10( T90 ),
       .io_in_9( T89 ),
       .io_in_8( T88 ),
       .io_in_7( T87 ),
       .io_in_6( T86 ),
       .io_in_5( T85 ),
       .io_in_4( T84 ),
       .io_in_3( T83 ),
       .io_in_2( T82 ),
       .io_in_1( T81 ),
       .io_in_0( T80 ),
       .io_out_15( streamMatrixTransposeTop_io_out_15 ),
       .io_out_14( streamMatrixTransposeTop_io_out_14 ),
       .io_out_13( streamMatrixTransposeTop_io_out_13 ),
       .io_out_12( streamMatrixTransposeTop_io_out_12 ),
       .io_out_11( streamMatrixTransposeTop_io_out_11 ),
       .io_out_10( streamMatrixTransposeTop_io_out_10 ),
       .io_out_9( streamMatrixTransposeTop_io_out_9 ),
       .io_out_8( streamMatrixTransposeTop_io_out_8 ),
       .io_out_7( streamMatrixTransposeTop_io_out_7 ),
       .io_out_6( streamMatrixTransposeTop_io_out_6 ),
       .io_out_5( streamMatrixTransposeTop_io_out_5 ),
       .io_out_4( streamMatrixTransposeTop_io_out_4 ),
       .io_out_3( streamMatrixTransposeTop_io_out_3 ),
       .io_out_2( streamMatrixTransposeTop_io_out_2 ),
       .io_out_1( streamMatrixTransposeTop_io_out_1 ),
       .io_out_0( streamMatrixTransposeTop_io_out_0 )
  );
  fft8_8 fft_2(.clk(clk), .reset(reset),
       .next( streamMatrixTransposeTop_io_start_next_stage ),
       .next_out( fft_2_next_out ),
       .X15( T79 ),
       .X14( T78 ),
       .X13( T77 ),
       .X12( T76 ),
       .X11( T75 ),
       .X10( T74 ),
       .X9( T73 ),
       .X8( T72 ),
       .X7( T71 ),
       .X6( T70 ),
       .X5( T69 ),
       .X4( T68 ),
       .X3( T67 ),
       .X2( T66 ),
       .X1( T65 ),
       .X0( T64 ),
       .Y15( fft_2_Y15 ),
       .Y14( fft_2_Y14 ),
       .Y13( fft_2_Y13 ),
       .Y12( fft_2_Y12 ),
       .Y11( fft_2_Y11 ),
       .Y10( fft_2_Y10 ),
       .Y9( fft_2_Y9 ),
       .Y8( fft_2_Y8 ),
       .Y7( fft_2_Y7 ),
       .Y6( fft_2_Y6 ),
       .Y5( fft_2_Y5 ),
       .Y4( fft_2_Y4 ),
       .Y3( fft_2_Y3 ),
       .Y2( fft_2_Y2 ),
       .Y1( fft_2_Y1 ),
       .Y0( fft_2_Y0 )
  );
  fft8_8 fft_3(.clk(clk), .reset(reset),
       .next( streamMatrixTransposeTop_io_start_next_stage ),
       //.next_out(  )
       .X15( T63 ),
       .X14( T62 ),
       .X13( T61 ),
       .X12( T60 ),
       .X11( T59 ),
       .X10( T58 ),
       .X9( T57 ),
       .X8( T56 ),
       .X7( T55 ),
       .X6( T54 ),
       .X5( T53 ),
       .X4( T52 ),
       .X3( T51 ),
       .X2( T50 ),
       .X1( T49 ),
       .X0( T48 ),
       .Y15( fft_3_Y15 ),
       .Y14( fft_3_Y14 ),
       .Y13( fft_3_Y13 ),
       .Y12( fft_3_Y12 ),
       .Y11( fft_3_Y11 ),
       .Y10( fft_3_Y10 ),
       .Y9( fft_3_Y9 ),
       .Y8( fft_3_Y8 ),
       .Y7( fft_3_Y7 ),
       .Y6( fft_3_Y6 ),
       .Y5( fft_3_Y5 ),
       .Y4( fft_3_Y4 ),
       .Y3( fft_3_Y3 ),
       .Y2( fft_3_Y2 ),
       .Y1( fft_3_Y1 ),
       .Y0( fft_3_Y0 )
  );
  multComplex multComplex(.clk(clk), .reset(reset),
       .io_real1( fft_2_Y0 ),
       .io_img1( fft_2_Y1 ),
       .io_real2( 32'h1 ),
       .io_img2( 32'h1 ),
       .io_realOut( multComplex_io_realOut ),
       .io_imgOut( multComplex_io_imgOut )
  );
  multComplex multComplex_1(.clk(clk), .reset(reset),
       .io_real1( fft_2_Y2 ),
       .io_img1( fft_2_Y3 ),
       .io_real2( 32'h1 ),
       .io_img2( 32'h1 ),
       .io_realOut( multComplex_1_io_realOut ),
       .io_imgOut( multComplex_1_io_imgOut )
  );
  multComplex multComplex_2(.clk(clk), .reset(reset),
       .io_real1( fft_2_Y4 ),
       .io_img1( fft_2_Y5 ),
       .io_real2( 32'h1 ),
       .io_img2( 32'h1 ),
       .io_realOut( multComplex_2_io_realOut ),
       .io_imgOut( multComplex_2_io_imgOut )
  );
  multComplex multComplex_3(.clk(clk), .reset(reset),
       .io_real1( fft_2_Y6 ),
       .io_img1( fft_2_Y7 ),
       .io_real2( 32'h1 ),
       .io_img2( 32'h1 ),
       .io_realOut( multComplex_3_io_realOut ),
       .io_imgOut( multComplex_3_io_imgOut )
  );
  multComplex multComplex_4(.clk(clk), .reset(reset),
       .io_real1( fft_2_Y8 ),
       .io_img1( fft_2_Y9 ),
       .io_real2( 32'h1 ),
       .io_img2( 32'h1 ),
       .io_realOut( multComplex_4_io_realOut ),
       .io_imgOut( multComplex_4_io_imgOut )
  );
  multComplex multComplex_5(.clk(clk), .reset(reset),
       .io_real1( fft_2_Y10 ),
       .io_img1( fft_2_Y11 ),
       .io_real2( 32'h1 ),
       .io_img2( 32'h1 ),
       .io_realOut( multComplex_5_io_realOut ),
       .io_imgOut( multComplex_5_io_imgOut )
  );
  multComplex multComplex_6(.clk(clk), .reset(reset),
       .io_real1( fft_2_Y12 ),
       .io_img1( fft_2_Y13 ),
       .io_real2( 32'h1 ),
       .io_img2( 32'h1 ),
       .io_realOut( multComplex_6_io_realOut ),
       .io_imgOut( multComplex_6_io_imgOut )
  );
  multComplex multComplex_7(.clk(clk), .reset(reset),
       .io_real1( fft_2_Y14 ),
       .io_img1( fft_2_Y15 ),
       .io_real2( 32'h1 ),
       .io_img2( 32'h1 ),
       .io_realOut( multComplex_7_io_realOut ),
       .io_imgOut( multComplex_7_io_imgOut )
  );
  multComplex multComplex_8(.clk(clk), .reset(reset),
       .io_real1( fft_3_Y0 ),
       .io_img1( fft_3_Y1 ),
       .io_real2( 32'h1 ),
       .io_img2( 32'h1 ),
       .io_realOut( multComplex_8_io_realOut ),
       .io_imgOut( multComplex_8_io_imgOut )
  );
  multComplex multComplex_9(.clk(clk), .reset(reset),
       .io_real1( fft_3_Y2 ),
       .io_img1( fft_3_Y3 ),
       .io_real2( 32'h1 ),
       .io_img2( 32'h1 ),
       .io_realOut( multComplex_9_io_realOut ),
       .io_imgOut( multComplex_9_io_imgOut )
  );
  multComplex multComplex_10(.clk(clk), .reset(reset),
       .io_real1( fft_3_Y4 ),
       .io_img1( fft_3_Y5 ),
       .io_real2( 32'h1 ),
       .io_img2( 32'h1 ),
       .io_realOut( multComplex_10_io_realOut ),
       .io_imgOut( multComplex_10_io_imgOut )
  );
  multComplex multComplex_11(.clk(clk), .reset(reset),
       .io_real1( fft_3_Y6 ),
       .io_img1( fft_3_Y7 ),
       .io_real2( 32'h1 ),
       .io_img2( 32'h1 ),
       .io_realOut( multComplex_11_io_realOut ),
       .io_imgOut( multComplex_11_io_imgOut )
  );
  multComplex multComplex_12(.clk(clk), .reset(reset),
       .io_real1( fft_3_Y8 ),
       .io_img1( fft_3_Y9 ),
       .io_real2( 32'h1 ),
       .io_img2( 32'h1 ),
       .io_realOut( multComplex_12_io_realOut ),
       .io_imgOut( multComplex_12_io_imgOut )
  );
  multComplex multComplex_13(.clk(clk), .reset(reset),
       .io_real1( fft_3_Y10 ),
       .io_img1( fft_3_Y11 ),
       .io_real2( 32'h1 ),
       .io_img2( 32'h1 ),
       .io_realOut( multComplex_13_io_realOut ),
       .io_imgOut( multComplex_13_io_imgOut )
  );
  multComplex multComplex_14(.clk(clk), .reset(reset),
       .io_real1( fft_3_Y12 ),
       .io_img1( fft_3_Y13 ),
       .io_real2( 32'h1 ),
       .io_img2( 32'h1 ),
       .io_realOut( multComplex_14_io_realOut ),
       .io_imgOut( multComplex_14_io_imgOut )
  );
  multComplex multComplex_15(.clk(clk), .reset(reset),
       .io_real1( fft_3_Y14 ),
       .io_img1( fft_3_Y15 ),
       .io_real2( 32'h1 ),
       .io_img2( 32'h1 ),
       .io_realOut( multComplex_15_io_realOut ),
       .io_imgOut( multComplex_15_io_imgOut )
  );
  ifft8_8 fft_4(.clk(clk), .reset(reset),
       .next( delayArrayNext_2 ),
       .next_out( fft_4_next_out ),
       .X15( multComplex_7_io_imgOut ),
       .X14( multComplex_7_io_realOut ),
       .X13( multComplex_6_io_imgOut ),
       .X12( multComplex_6_io_realOut ),
       .X11( multComplex_5_io_imgOut ),
       .X10( multComplex_5_io_realOut ),
       .X9( multComplex_4_io_imgOut ),
       .X8( multComplex_4_io_realOut ),
       .X7( multComplex_3_io_imgOut ),
       .X6( multComplex_3_io_realOut ),
       .X5( multComplex_2_io_imgOut ),
       .X4( multComplex_2_io_realOut ),
       .X3( multComplex_1_io_imgOut ),
       .X2( multComplex_1_io_realOut ),
       .X1( multComplex_io_imgOut ),
       .X0( multComplex_io_realOut ),
       .Y15( fft_4_Y15 ),
       .Y14( fft_4_Y14 ),
       .Y13( fft_4_Y13 ),
       .Y12( fft_4_Y12 ),
       .Y11( fft_4_Y11 ),
       .Y10( fft_4_Y10 ),
       .Y9( fft_4_Y9 ),
       .Y8( fft_4_Y8 ),
       .Y7( fft_4_Y7 ),
       .Y6( fft_4_Y6 ),
       .Y5( fft_4_Y5 ),
       .Y4( fft_4_Y4 ),
       .Y3( fft_4_Y3 ),
       .Y2( fft_4_Y2 ),
       .Y1( fft_4_Y1 ),
       .Y0( fft_4_Y0 )
  );
  ifft8_8 fft_5(.clk(clk), .reset(reset),
       .next( delayArrayNext_2 ),
       //.next_out(  )
       .X15( multComplex_15_io_imgOut ),
       .X14( multComplex_15_io_realOut ),
       .X13( multComplex_14_io_imgOut ),
       .X12( multComplex_14_io_realOut ),
       .X11( multComplex_13_io_imgOut ),
       .X10( multComplex_13_io_realOut ),
       .X9( multComplex_12_io_imgOut ),
       .X8( multComplex_12_io_realOut ),
       .X7( multComplex_11_io_imgOut ),
       .X6( multComplex_11_io_realOut ),
       .X5( multComplex_10_io_imgOut ),
       .X4( multComplex_10_io_realOut ),
       .X3( multComplex_9_io_imgOut ),
       .X2( multComplex_9_io_realOut ),
       .X1( multComplex_8_io_imgOut ),
       .X0( multComplex_8_io_realOut ),
       .Y15( fft_5_Y15 ),
       .Y14( fft_5_Y14 ),
       .Y13( fft_5_Y13 ),
       .Y12( fft_5_Y12 ),
       .Y11( fft_5_Y11 ),
       .Y10( fft_5_Y10 ),
       .Y9( fft_5_Y9 ),
       .Y8( fft_5_Y8 ),
       .Y7( fft_5_Y7 ),
       .Y6( fft_5_Y6 ),
       .Y5( fft_5_Y5 ),
       .Y4( fft_5_Y4 ),
       .Y3( fft_5_Y3 ),
       .Y2( fft_5_Y2 ),
       .Y1( fft_5_Y1 ),
       .Y0( fft_5_Y0 )
  );
  ifft8_8 fft_6(.clk(clk), .reset(reset),
       .next( streamMatrixTransposeTop_1_io_start_next_stage ),
       .next_out( fft_6_next_out ),
       .X15( T47 ),
       .X14( T46 ),
       .X13( T45 ),
       .X12( T44 ),
       .X11( T43 ),
       .X10( T42 ),
       .X9( T41 ),
       .X8( T40 ),
       .X7( T39 ),
       .X6( T38 ),
       .X5( T37 ),
       .X4( T36 ),
       .X3( T35 ),
       .X2( T34 ),
       .X1( T33 ),
       .X0( T32 ),
       //.Y15(  )
       .Y14( fft_6_Y14 ),
       //.Y13(  )
       .Y12( fft_6_Y12 ),
       //.Y11(  )
       .Y10( fft_6_Y10 ),
       //.Y9(  )
       .Y8( fft_6_Y8 ),
       //.Y7(  )
       .Y6( fft_6_Y6 ),
       //.Y5(  )
       .Y4( fft_6_Y4 ),
       //.Y3(  )
       .Y2( fft_6_Y2 ),
       //.Y1(  )
       .Y0( fft_6_Y0 )
  );
  ifft8_8 fft_7(.clk(clk), .reset(reset),
       .next( streamMatrixTransposeTop_1_io_start_next_stage ),
       //.next_out(  )
       .X15( T31 ),
       .X14( T30 ),
       .X13( T29 ),
       .X12( T28 ),
       .X11( T27 ),
       .X10( T26 ),
       .X9( T25 ),
       .X8( T24 ),
       .X7( T23 ),
       .X6( T22 ),
       .X5( T21 ),
       .X4( T20 ),
       .X3( T19 ),
       .X2( T18 ),
       .X1( T17 ),
       .X0( T16 ),
       //.Y15(  )
       .Y14( fft_7_Y14 ),
       //.Y13(  )
       .Y12( fft_7_Y12 ),
       //.Y11(  )
       .Y10( fft_7_Y10 ),
       //.Y9(  )
       .Y8( fft_7_Y8 ),
       //.Y7(  )
       .Y6( fft_7_Y6 ),
       //.Y5(  )
       .Y4( fft_7_Y4 ),
       //.Y3(  )
       .Y2( fft_7_Y2 ),
       //.Y1(  )
       .Y0( fft_7_Y0 )
  );
  streamMatrixTransposeTop streamMatrixTransposeTop_1(.clk(clk), .reset(reset),
       .io_clk_en( 1'h1 ),
       .io_start( startSecondMatrix ),
       .io_start_next_stage( streamMatrixTransposeTop_1_io_start_next_stage ),
       .io_in_15( T15 ),
       .io_in_14( T14 ),
       .io_in_13( T13 ),
       .io_in_12( T12 ),
       .io_in_11( T11 ),
       .io_in_10( T10 ),
       .io_in_9( T9 ),
       .io_in_8( T8 ),
       .io_in_7( T7 ),
       .io_in_6( T6 ),
       .io_in_5( T5 ),
       .io_in_4( T4 ),
       .io_in_3( T3 ),
       .io_in_2( T2 ),
       .io_in_1( T1 ),
       .io_in_0( T0 ),
       .io_out_15( streamMatrixTransposeTop_1_io_out_15 ),
       .io_out_14( streamMatrixTransposeTop_1_io_out_14 ),
       .io_out_13( streamMatrixTransposeTop_1_io_out_13 ),
       .io_out_12( streamMatrixTransposeTop_1_io_out_12 ),
       .io_out_11( streamMatrixTransposeTop_1_io_out_11 ),
       .io_out_10( streamMatrixTransposeTop_1_io_out_10 ),
       .io_out_9( streamMatrixTransposeTop_1_io_out_9 ),
       .io_out_8( streamMatrixTransposeTop_1_io_out_8 ),
       .io_out_7( streamMatrixTransposeTop_1_io_out_7 ),
       .io_out_6( streamMatrixTransposeTop_1_io_out_6 ),
       .io_out_5( streamMatrixTransposeTop_1_io_out_5 ),
       .io_out_4( streamMatrixTransposeTop_1_io_out_4 ),
       .io_out_3( streamMatrixTransposeTop_1_io_out_3 ),
       .io_out_2( streamMatrixTransposeTop_1_io_out_2 ),
       .io_out_1( streamMatrixTransposeTop_1_io_out_1 ),
       .io_out_0( streamMatrixTransposeTop_1_io_out_0 )
  );

  always @(posedge clk) begin
    startSecondMatrix <= fft_4_next_out;
    delaySecond_8 <= streamMatrixTransposeTop_1_io_out_8;
    delaySecond_9 <= streamMatrixTransposeTop_1_io_out_9;
    delaySecond_10 <= streamMatrixTransposeTop_1_io_out_10;
    delaySecond_11 <= streamMatrixTransposeTop_1_io_out_11;
    delaySecond_12 <= streamMatrixTransposeTop_1_io_out_12;
    delaySecond_13 <= streamMatrixTransposeTop_1_io_out_13;
    delaySecond_14 <= streamMatrixTransposeTop_1_io_out_14;
    delaySecond_15 <= streamMatrixTransposeTop_1_io_out_15;
    delaySecond_0 <= streamMatrixTransposeTop_1_io_out_0;
    delaySecond_1 <= streamMatrixTransposeTop_1_io_out_1;
    delaySecond_2 <= streamMatrixTransposeTop_1_io_out_2;
    delaySecond_3 <= streamMatrixTransposeTop_1_io_out_3;
    delaySecond_4 <= streamMatrixTransposeTop_1_io_out_4;
    delaySecond_5 <= streamMatrixTransposeTop_1_io_out_5;
    delaySecond_6 <= streamMatrixTransposeTop_1_io_out_6;
    delaySecond_7 <= streamMatrixTransposeTop_1_io_out_7;
    delayArrayNext_2 <= delayArrayNext_1;
    delayArrayNext_1 <= delayArrayNext_0;
    delayArrayNext_0 <= fft_2_next_out;
    delayFirst_8 <= streamMatrixTransposeTop_io_out_8;
    delayFirst_9 <= streamMatrixTransposeTop_io_out_9;
    delayFirst_10 <= streamMatrixTransposeTop_io_out_10;
    delayFirst_11 <= streamMatrixTransposeTop_io_out_11;
    delayFirst_12 <= streamMatrixTransposeTop_io_out_12;
    delayFirst_13 <= streamMatrixTransposeTop_io_out_13;
    delayFirst_14 <= streamMatrixTransposeTop_io_out_14;
    delayFirst_15 <= streamMatrixTransposeTop_io_out_15;
    delayFirst_0 <= streamMatrixTransposeTop_io_out_0;
    delayFirst_1 <= streamMatrixTransposeTop_io_out_1;
    delayFirst_2 <= streamMatrixTransposeTop_io_out_2;
    delayFirst_3 <= streamMatrixTransposeTop_io_out_3;
    delayFirst_4 <= streamMatrixTransposeTop_io_out_4;
    delayFirst_5 <= streamMatrixTransposeTop_io_out_5;
    delayFirst_6 <= streamMatrixTransposeTop_io_out_6;
    delayFirst_7 <= streamMatrixTransposeTop_io_out_7;
    startFirstMatrix <= fft_next_out;
    delayInput_8 <= io_in_8;
    delayInput_9 <= io_in_9;
    delayInput_10 <= io_in_10;
    delayInput_11 <= io_in_11;
    delayInput_12 <= io_in_12;
    delayInput_13 <= io_in_13;
    delayInput_14 <= io_in_14;
    delayInput_15 <= io_in_15;
    delayInput_0 <= io_in_0;
    delayInput_1 <= io_in_1;
    delayInput_2 <= io_in_2;
    delayInput_3 <= io_in_3;
    delayInput_4 <= io_in_4;
    delayInput_5 <= io_in_5;
    delayInput_6 <= io_in_6;
    delayInput_7 <= io_in_7;
    delayStartNextStage <= fft_6_next_out;
  end
endmodule

module afu_user(input clk, input reset,
    input [511:0] input_fifo_din,
    input  input_fifo_we,
    output input_fifo_full,
    output input_fifo_almost_full,
    output[5:0] input_fifo_count,
    output[511:0] output_fifo_dout,
    input  output_fifo_re,
    output output_fifo_empty,
    output output_fifo_almost_empty,
    input [31:0] ctx_length
);

  wire T0;
  wire T1;
  wire T2;
  reg [31:0] ctx_output_count;
  wire[31:0] T46;
  wire[31:0] T3;
  wire[31:0] T4;
  wire[511:0] T5;
  wire[511:0] T6;
  wire[255:0] T7;
  wire[127:0] T8;
  wire[63:0] T9;
  wire[63:0] T10;
  wire[127:0] T11;
  wire[63:0] T12;
  wire[63:0] T13;
  wire[255:0] T14;
  wire[127:0] T15;
  wire[63:0] T16;
  wire[63:0] T17;
  wire[127:0] T18;
  wire[63:0] T19;
  wire[63:0] T20;
  wire[31:0] T21;
  wire[31:0] T22;
  wire[31:0] T23;
  wire[31:0] T24;
  wire[31:0] T25;
  wire[31:0] T26;
  wire[31:0] T27;
  wire[31:0] T28;
  wire[31:0] T29;
  wire[31:0] T30;
  wire[31:0] T31;
  wire[31:0] T32;
  wire[31:0] T33;
  wire[31:0] T34;
  wire[31:0] T35;
  wire[31:0] T36;
  reg  start_reg;
  wire T47;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  reg [31:0] ctx_input_count;
  wire[31:0] T48;
  wire[31:0] T42;
  wire[31:0] T43;
  wire T44;
  wire T45;
  wire[5:0] T49;
  wire[511:0] syn_read_fifo_dout;
  wire syn_read_fifo_empty;
  wire syn_read_fifo_full;
  wire syn_read_fifo_count;
  wire syn_read_fifo_almostfull;
  wire[511:0] syn_read_fifo_1_dout;
  wire syn_read_fifo_1_empty;
  wire syn_read_fifo_1_almostempty;
  wire two_d_convolution_io_start_next_stage;
  wire[31:0] two_d_convolution_io_out_15;
  wire[31:0] two_d_convolution_io_out_14;
  wire[31:0] two_d_convolution_io_out_13;
  wire[31:0] two_d_convolution_io_out_12;
  wire[31:0] two_d_convolution_io_out_11;
  wire[31:0] two_d_convolution_io_out_10;
  wire[31:0] two_d_convolution_io_out_9;
  wire[31:0] two_d_convolution_io_out_8;
  wire[31:0] two_d_convolution_io_out_7;
  wire[31:0] two_d_convolution_io_out_6;
  wire[31:0] two_d_convolution_io_out_5;
  wire[31:0] two_d_convolution_io_out_4;
  wire[31:0] two_d_convolution_io_out_3;
  wire[31:0] two_d_convolution_io_out_2;
  wire[31:0] two_d_convolution_io_out_1;
  wire[31:0] two_d_convolution_io_out_0;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    ctx_output_count = {1{$random}};
    start_reg = {1{$random}};
    ctx_input_count = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = T2 ? 1'h0 : T1;
  assign T1 = two_d_convolution_io_start_next_stage & T40;
  assign T2 = ctx_length == ctx_output_count;
  assign T46 = reset ? 32'h0 : T3;
  assign T3 = T0 ? T4 : ctx_output_count;
  assign T4 = ctx_output_count + 32'h1;
  assign T5 = T6;
  assign T6 = {T14, T7};
  assign T7 = {T11, T8};
  assign T8 = {T10, T9};
  assign T9 = {two_d_convolution_io_out_1, two_d_convolution_io_out_0};
  assign T10 = {two_d_convolution_io_out_3, two_d_convolution_io_out_2};
  assign T11 = {T13, T12};
  assign T12 = {two_d_convolution_io_out_5, two_d_convolution_io_out_4};
  assign T13 = {two_d_convolution_io_out_7, two_d_convolution_io_out_6};
  assign T14 = {T18, T15};
  assign T15 = {T17, T16};
  assign T16 = {two_d_convolution_io_out_9, two_d_convolution_io_out_8};
  assign T17 = {two_d_convolution_io_out_11, two_d_convolution_io_out_10};
  assign T18 = {T20, T19};
  assign T19 = {two_d_convolution_io_out_13, two_d_convolution_io_out_12};
  assign T20 = {two_d_convolution_io_out_15, two_d_convolution_io_out_14};
  assign T21 = syn_read_fifo_dout[31:0];
  assign T22 = syn_read_fifo_dout[63:32];
  assign T23 = syn_read_fifo_dout[95:64];
  assign T24 = syn_read_fifo_dout[127:96];
  assign T25 = syn_read_fifo_dout[159:128];
  assign T26 = syn_read_fifo_dout[191:160];
  assign T27 = syn_read_fifo_dout[223:192];
  assign T28 = syn_read_fifo_dout[255:224];
  assign T29 = syn_read_fifo_dout[287:256];
  assign T30 = syn_read_fifo_dout[319:288];
  assign T31 = syn_read_fifo_dout[351:320];
  assign T32 = syn_read_fifo_dout[383:352];
  assign T33 = syn_read_fifo_dout[415:384];
  assign T34 = syn_read_fifo_dout[447:416];
  assign T35 = syn_read_fifo_dout[479:448];
  assign T36 = syn_read_fifo_dout[511:480];
  assign T47 = reset ? 1'h0 : T37;
  assign T37 = T39 ? 1'h0 : T38;
  assign T38 = T44 ? 1'h1 : start_reg;
  assign T39 = T44 ^ 1'h1;
  assign T40 = T41 ? 1'h1 : start_reg;
  assign T41 = ctx_length == ctx_input_count;
  assign T48 = reset ? 32'h0 : T42;
  assign T42 = T44 ? T43 : ctx_input_count;
  assign T43 = ctx_input_count + 32'h1;
  assign T44 = reset ? 1'h0 : T45;
  assign T45 = ~ syn_read_fifo_empty;
  assign output_fifo_almost_empty = syn_read_fifo_1_almostempty;
  assign output_fifo_empty = syn_read_fifo_1_empty;
  assign output_fifo_dout = syn_read_fifo_1_dout;
  assign input_fifo_count = T49;
  assign T49 = {5'h0, syn_read_fifo_count};
  assign input_fifo_almost_full = syn_read_fifo_almostfull;
  assign input_fifo_full = syn_read_fifo_full;
  syn_read_fifo #(.FIFO_WIDTH(512),.FIFO_DEPTH_BITS(6),.FIFO_ALMOSTFULL_THRESHOLD(60),.FIFO_ALMOSTEMPTY_THRESHOLD(2))
  syn_read_fifo(.clk(clk), .reset(reset),
       .din( input_fifo_din ),
       .we( input_fifo_we ),
       .re( T44 ),
       .dout( syn_read_fifo_dout ),
       .empty( syn_read_fifo_empty ),
       //.almostempty(  )
       .full( syn_read_fifo_full ),
       .count( syn_read_fifo_count ),
       .almostfull( syn_read_fifo_almostfull )
  );
  two_d_convolution two_d_convolution(.clk(clk), .reset(reset),
       .io_clk_en( T40 ),
       .io_start( start_reg ),
       .io_start_next_stage( two_d_convolution_io_start_next_stage ),
       .io_in_15( T36 ),
       .io_in_14( T35 ),
       .io_in_13( T34 ),
       .io_in_12( T33 ),
       .io_in_11( T32 ),
       .io_in_10( T31 ),
       .io_in_9( T30 ),
       .io_in_8( T29 ),
       .io_in_7( T28 ),
       .io_in_6( T27 ),
       .io_in_5( T26 ),
       .io_in_4( T25 ),
       .io_in_3( T24 ),
       .io_in_2( T23 ),
       .io_in_1( T22 ),
       .io_in_0( T21 ),
       .io_out_15( two_d_convolution_io_out_15 ),
       .io_out_14( two_d_convolution_io_out_14 ),
       .io_out_13( two_d_convolution_io_out_13 ),
       .io_out_12( two_d_convolution_io_out_12 ),
       .io_out_11( two_d_convolution_io_out_11 ),
       .io_out_10( two_d_convolution_io_out_10 ),
       .io_out_9( two_d_convolution_io_out_9 ),
       .io_out_8( two_d_convolution_io_out_8 ),
       .io_out_7( two_d_convolution_io_out_7 ),
       .io_out_6( two_d_convolution_io_out_6 ),
       .io_out_5( two_d_convolution_io_out_5 ),
       .io_out_4( two_d_convolution_io_out_4 ),
       .io_out_3( two_d_convolution_io_out_3 ),
       .io_out_2( two_d_convolution_io_out_2 ),
       .io_out_1( two_d_convolution_io_out_1 ),
       .io_out_0( two_d_convolution_io_out_0 )
  );
  syn_read_fifo #(.FIFO_WIDTH(512),.FIFO_DEPTH_BITS(6),.FIFO_ALMOSTFULL_THRESHOLD(60),.FIFO_ALMOSTEMPTY_THRESHOLD(2))
  syn_read_fifo_1(.clk(clk), .reset(reset),
       .din( T5 ),
       .we( T0 ),
       .re( output_fifo_re ),
       .dout( syn_read_fifo_1_dout ),
       .empty( syn_read_fifo_1_empty ),
       .almostempty( syn_read_fifo_1_almostempty )
       //.full(  )
       //.count(  )
       //.almostfull(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      ctx_output_count <= 32'h0;
    end else if(T0) begin
      ctx_output_count <= T4;
    end
    if(reset) begin
      start_reg <= 1'h0;
    end else if(T39) begin
      start_reg <= 1'h0;
    end else if(T44) begin
      start_reg <= 1'h1;
    end
    if(reset) begin
      ctx_input_count <= 32'h0;
    end else if(T44) begin
      ctx_input_count <= T43;
    end
  end
endmodule

