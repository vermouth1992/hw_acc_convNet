module crossbar(input clk, input reset,
    input  io_clk_en,
    input  io_start,
    output io_start_next_stage,
    input [31:0] io_in_31,
    input [31:0] io_in_30,
    input [31:0] io_in_29,
    input [31:0] io_in_28,
    input [31:0] io_in_27,
    input [31:0] io_in_26,
    input [31:0] io_in_25,
    input [31:0] io_in_24,
    input [31:0] io_in_23,
    input [31:0] io_in_22,
    input [31:0] io_in_21,
    input [31:0] io_in_20,
    input [31:0] io_in_19,
    input [31:0] io_in_18,
    input [31:0] io_in_17,
    input [31:0] io_in_16,
    input [31:0] io_in_15,
    input [31:0] io_in_14,
    input [31:0] io_in_13,
    input [31:0] io_in_12,
    input [31:0] io_in_11,
    input [31:0] io_in_10,
    input [31:0] io_in_9,
    input [31:0] io_in_8,
    input [31:0] io_in_7,
    input [31:0] io_in_6,
    input [31:0] io_in_5,
    input [31:0] io_in_4,
    input [31:0] io_in_3,
    input [31:0] io_in_2,
    input [31:0] io_in_1,
    input [31:0] io_in_0,
    output[31:0] io_out_31,
    output[31:0] io_out_30,
    output[31:0] io_out_29,
    output[31:0] io_out_28,
    output[31:0] io_out_27,
    output[31:0] io_out_26,
    output[31:0] io_out_25,
    output[31:0] io_out_24,
    output[31:0] io_out_23,
    output[31:0] io_out_22,
    output[31:0] io_out_21,
    output[31:0] io_out_20,
    output[31:0] io_out_19,
    output[31:0] io_out_18,
    output[31:0] io_out_17,
    output[31:0] io_out_16,
    output[31:0] io_out_15,
    output[31:0] io_out_14,
    output[31:0] io_out_13,
    output[31:0] io_out_12,
    output[31:0] io_out_11,
    output[31:0] io_out_10,
    output[31:0] io_out_9,
    output[31:0] io_out_8,
    output[31:0] io_out_7,
    output[31:0] io_out_6,
    output[31:0] io_out_5,
    output[31:0] io_out_4,
    output[31:0] io_out_3,
    output[31:0] io_out_2,
    output[31:0] io_out_1,
    output[31:0] io_out_0
);

  reg [31:0] out_reg_0;
  wire[31:0] T0;
  wire T1;
  reg [31:0] out_reg_1;
  wire[31:0] T2;
  reg [31:0] out_reg_2;
  wire[31:0] T3;
  reg [31:0] out_reg_3;
  wire[31:0] T4;
  reg [31:0] out_reg_4;
  wire[31:0] T5;
  reg [31:0] out_reg_5;
  wire[31:0] T6;
  reg [31:0] out_reg_6;
  wire[31:0] T7;
  reg [31:0] out_reg_7;
  wire[31:0] T8;
  reg [31:0] out_reg_8;
  wire[31:0] T9;
  reg [31:0] out_reg_9;
  wire[31:0] T10;
  reg [31:0] out_reg_10;
  wire[31:0] T11;
  reg [31:0] out_reg_11;
  wire[31:0] T12;
  reg [31:0] out_reg_12;
  wire[31:0] T13;
  reg [31:0] out_reg_13;
  wire[31:0] T14;
  reg [31:0] out_reg_14;
  wire[31:0] T15;
  reg [31:0] out_reg_15;
  wire[31:0] T16;
  reg [31:0] out_reg_16;
  wire[31:0] T17;
  reg [31:0] out_reg_17;
  wire[31:0] T18;
  reg [31:0] out_reg_18;
  wire[31:0] T19;
  reg [31:0] out_reg_19;
  wire[31:0] T20;
  reg [31:0] out_reg_20;
  wire[31:0] T21;
  reg [31:0] out_reg_21;
  wire[31:0] T22;
  reg [31:0] out_reg_22;
  wire[31:0] T23;
  reg [31:0] out_reg_23;
  wire[31:0] T24;
  reg [31:0] out_reg_24;
  wire[31:0] T25;
  reg [31:0] out_reg_25;
  wire[31:0] T26;
  reg [31:0] out_reg_26;
  wire[31:0] T27;
  reg [31:0] out_reg_27;
  wire[31:0] T28;
  reg [31:0] out_reg_28;
  wire[31:0] T29;
  reg [31:0] out_reg_29;
  wire[31:0] T30;
  reg [31:0] out_reg_30;
  wire[31:0] T31;
  reg [31:0] out_reg_31;
  wire[31:0] T32;
  reg  start_next_stage_reg;
  wire T35;
  wire T33;
  wire T34;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    out_reg_0 = {1{$random}};
    out_reg_1 = {1{$random}};
    out_reg_2 = {1{$random}};
    out_reg_3 = {1{$random}};
    out_reg_4 = {1{$random}};
    out_reg_5 = {1{$random}};
    out_reg_6 = {1{$random}};
    out_reg_7 = {1{$random}};
    out_reg_8 = {1{$random}};
    out_reg_9 = {1{$random}};
    out_reg_10 = {1{$random}};
    out_reg_11 = {1{$random}};
    out_reg_12 = {1{$random}};
    out_reg_13 = {1{$random}};
    out_reg_14 = {1{$random}};
    out_reg_15 = {1{$random}};
    out_reg_16 = {1{$random}};
    out_reg_17 = {1{$random}};
    out_reg_18 = {1{$random}};
    out_reg_19 = {1{$random}};
    out_reg_20 = {1{$random}};
    out_reg_21 = {1{$random}};
    out_reg_22 = {1{$random}};
    out_reg_23 = {1{$random}};
    out_reg_24 = {1{$random}};
    out_reg_25 = {1{$random}};
    out_reg_26 = {1{$random}};
    out_reg_27 = {1{$random}};
    out_reg_28 = {1{$random}};
    out_reg_29 = {1{$random}};
    out_reg_30 = {1{$random}};
    out_reg_31 = {1{$random}};
    start_next_stage_reg = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_out_0 = out_reg_0;
  assign T0 = T1 ? io_in_0 : out_reg_0;
  assign T1 = io_clk_en & io_start;
  assign io_out_1 = out_reg_1;
  assign T2 = T1 ? io_in_8 : out_reg_1;
  assign io_out_2 = out_reg_2;
  assign T3 = T1 ? io_in_16 : out_reg_2;
  assign io_out_3 = out_reg_3;
  assign T4 = T1 ? io_in_24 : out_reg_3;
  assign io_out_4 = out_reg_4;
  assign T5 = T1 ? io_in_4 : out_reg_4;
  assign io_out_5 = out_reg_5;
  assign T6 = T1 ? io_in_12 : out_reg_5;
  assign io_out_6 = out_reg_6;
  assign T7 = T1 ? io_in_20 : out_reg_6;
  assign io_out_7 = out_reg_7;
  assign T8 = T1 ? io_in_28 : out_reg_7;
  assign io_out_8 = out_reg_8;
  assign T9 = T1 ? io_in_1 : out_reg_8;
  assign io_out_9 = out_reg_9;
  assign T10 = T1 ? io_in_9 : out_reg_9;
  assign io_out_10 = out_reg_10;
  assign T11 = T1 ? io_in_17 : out_reg_10;
  assign io_out_11 = out_reg_11;
  assign T12 = T1 ? io_in_25 : out_reg_11;
  assign io_out_12 = out_reg_12;
  assign T13 = T1 ? io_in_5 : out_reg_12;
  assign io_out_13 = out_reg_13;
  assign T14 = T1 ? io_in_13 : out_reg_13;
  assign io_out_14 = out_reg_14;
  assign T15 = T1 ? io_in_21 : out_reg_14;
  assign io_out_15 = out_reg_15;
  assign T16 = T1 ? io_in_29 : out_reg_15;
  assign io_out_16 = out_reg_16;
  assign T17 = T1 ? io_in_2 : out_reg_16;
  assign io_out_17 = out_reg_17;
  assign T18 = T1 ? io_in_10 : out_reg_17;
  assign io_out_18 = out_reg_18;
  assign T19 = T1 ? io_in_18 : out_reg_18;
  assign io_out_19 = out_reg_19;
  assign T20 = T1 ? io_in_26 : out_reg_19;
  assign io_out_20 = out_reg_20;
  assign T21 = T1 ? io_in_6 : out_reg_20;
  assign io_out_21 = out_reg_21;
  assign T22 = T1 ? io_in_14 : out_reg_21;
  assign io_out_22 = out_reg_22;
  assign T23 = T1 ? io_in_22 : out_reg_22;
  assign io_out_23 = out_reg_23;
  assign T24 = T1 ? io_in_30 : out_reg_23;
  assign io_out_24 = out_reg_24;
  assign T25 = T1 ? io_in_3 : out_reg_24;
  assign io_out_25 = out_reg_25;
  assign T26 = T1 ? io_in_11 : out_reg_25;
  assign io_out_26 = out_reg_26;
  assign T27 = T1 ? io_in_19 : out_reg_26;
  assign io_out_27 = out_reg_27;
  assign T28 = T1 ? io_in_27 : out_reg_27;
  assign io_out_28 = out_reg_28;
  assign T29 = T1 ? io_in_7 : out_reg_28;
  assign io_out_29 = out_reg_29;
  assign T30 = T1 ? io_in_15 : out_reg_29;
  assign io_out_30 = out_reg_30;
  assign T31 = T1 ? io_in_23 : out_reg_30;
  assign io_out_31 = out_reg_31;
  assign T32 = T1 ? io_in_31 : out_reg_31;
  assign io_start_next_stage = start_next_stage_reg;
  assign T35 = reset ? 1'h0 : T33;
  assign T33 = T34 ? 1'h1 : start_next_stage_reg;
  assign T34 = io_start & io_clk_en;

  always @(posedge clk) begin
    if(T1) begin
      out_reg_0 <= io_in_0;
    end
    if(T1) begin
      out_reg_1 <= io_in_8;
    end
    if(T1) begin
      out_reg_2 <= io_in_16;
    end
    if(T1) begin
      out_reg_3 <= io_in_24;
    end
    if(T1) begin
      out_reg_4 <= io_in_4;
    end
    if(T1) begin
      out_reg_5 <= io_in_12;
    end
    if(T1) begin
      out_reg_6 <= io_in_20;
    end
    if(T1) begin
      out_reg_7 <= io_in_28;
    end
    if(T1) begin
      out_reg_8 <= io_in_1;
    end
    if(T1) begin
      out_reg_9 <= io_in_9;
    end
    if(T1) begin
      out_reg_10 <= io_in_17;
    end
    if(T1) begin
      out_reg_11 <= io_in_25;
    end
    if(T1) begin
      out_reg_12 <= io_in_5;
    end
    if(T1) begin
      out_reg_13 <= io_in_13;
    end
    if(T1) begin
      out_reg_14 <= io_in_21;
    end
    if(T1) begin
      out_reg_15 <= io_in_29;
    end
    if(T1) begin
      out_reg_16 <= io_in_2;
    end
    if(T1) begin
      out_reg_17 <= io_in_10;
    end
    if(T1) begin
      out_reg_18 <= io_in_18;
    end
    if(T1) begin
      out_reg_19 <= io_in_26;
    end
    if(T1) begin
      out_reg_20 <= io_in_6;
    end
    if(T1) begin
      out_reg_21 <= io_in_14;
    end
    if(T1) begin
      out_reg_22 <= io_in_22;
    end
    if(T1) begin
      out_reg_23 <= io_in_30;
    end
    if(T1) begin
      out_reg_24 <= io_in_3;
    end
    if(T1) begin
      out_reg_25 <= io_in_11;
    end
    if(T1) begin
      out_reg_26 <= io_in_19;
    end
    if(T1) begin
      out_reg_27 <= io_in_27;
    end
    if(T1) begin
      out_reg_28 <= io_in_7;
    end
    if(T1) begin
      out_reg_29 <= io_in_15;
    end
    if(T1) begin
      out_reg_30 <= io_in_23;
    end
    if(T1) begin
      out_reg_31 <= io_in_31;
    end
    if(reset) begin
      start_next_stage_reg <= 1'h0;
    end else if(T34) begin
      start_next_stage_reg <= 1'h1;
    end
  end
endmodule

module crossbarShiftDown(input clk, input reset,
    input  io_clk_en,
    input  io_start,
    output io_start_next_stage,
    input [31:0] io_in_31,
    input [31:0] io_in_30,
    input [31:0] io_in_29,
    input [31:0] io_in_28,
    input [31:0] io_in_27,
    input [31:0] io_in_26,
    input [31:0] io_in_25,
    input [31:0] io_in_24,
    input [31:0] io_in_23,
    input [31:0] io_in_22,
    input [31:0] io_in_21,
    input [31:0] io_in_20,
    input [31:0] io_in_19,
    input [31:0] io_in_18,
    input [31:0] io_in_17,
    input [31:0] io_in_16,
    input [31:0] io_in_15,
    input [31:0] io_in_14,
    input [31:0] io_in_13,
    input [31:0] io_in_12,
    input [31:0] io_in_11,
    input [31:0] io_in_10,
    input [31:0] io_in_9,
    input [31:0] io_in_8,
    input [31:0] io_in_7,
    input [31:0] io_in_6,
    input [31:0] io_in_5,
    input [31:0] io_in_4,
    input [31:0] io_in_3,
    input [31:0] io_in_2,
    input [31:0] io_in_1,
    input [31:0] io_in_0,
    output[31:0] io_out_31,
    output[31:0] io_out_30,
    output[31:0] io_out_29,
    output[31:0] io_out_28,
    output[31:0] io_out_27,
    output[31:0] io_out_26,
    output[31:0] io_out_25,
    output[31:0] io_out_24,
    output[31:0] io_out_23,
    output[31:0] io_out_22,
    output[31:0] io_out_21,
    output[31:0] io_out_20,
    output[31:0] io_out_19,
    output[31:0] io_out_18,
    output[31:0] io_out_17,
    output[31:0] io_out_16,
    output[31:0] io_out_15,
    output[31:0] io_out_14,
    output[31:0] io_out_13,
    output[31:0] io_out_12,
    output[31:0] io_out_11,
    output[31:0] io_out_10,
    output[31:0] io_out_9,
    output[31:0] io_out_8,
    output[31:0] io_out_7,
    output[31:0] io_out_6,
    output[31:0] io_out_5,
    output[31:0] io_out_4,
    output[31:0] io_out_3,
    output[31:0] io_out_2,
    output[31:0] io_out_1,
    output[31:0] io_out_0
);

  reg [31:0] out_reg_0;
  wire[31:0] T0;
  wire[31:0] T1;
  wire T2;
  wire T3;
  reg  timestamp;
  wire T73;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  reg [31:0] out_reg_1;
  wire[31:0] T10;
  wire[31:0] T11;
  reg [31:0] out_reg_2;
  wire[31:0] T12;
  wire[31:0] T13;
  reg [31:0] out_reg_3;
  wire[31:0] T14;
  wire[31:0] T15;
  reg [31:0] out_reg_4;
  wire[31:0] T16;
  wire[31:0] T17;
  reg [31:0] out_reg_5;
  wire[31:0] T18;
  wire[31:0] T19;
  reg [31:0] out_reg_6;
  wire[31:0] T20;
  wire[31:0] T21;
  reg [31:0] out_reg_7;
  wire[31:0] T22;
  wire[31:0] T23;
  reg [31:0] out_reg_8;
  wire[31:0] T24;
  wire[31:0] T25;
  reg [31:0] out_reg_9;
  wire[31:0] T26;
  wire[31:0] T27;
  reg [31:0] out_reg_10;
  wire[31:0] T28;
  wire[31:0] T29;
  reg [31:0] out_reg_11;
  wire[31:0] T30;
  wire[31:0] T31;
  reg [31:0] out_reg_12;
  wire[31:0] T32;
  wire[31:0] T33;
  reg [31:0] out_reg_13;
  wire[31:0] T34;
  wire[31:0] T35;
  reg [31:0] out_reg_14;
  wire[31:0] T36;
  wire[31:0] T37;
  reg [31:0] out_reg_15;
  wire[31:0] T38;
  wire[31:0] T39;
  reg [31:0] out_reg_16;
  wire[31:0] T40;
  wire[31:0] T41;
  reg [31:0] out_reg_17;
  wire[31:0] T42;
  wire[31:0] T43;
  reg [31:0] out_reg_18;
  wire[31:0] T44;
  wire[31:0] T45;
  reg [31:0] out_reg_19;
  wire[31:0] T46;
  wire[31:0] T47;
  reg [31:0] out_reg_20;
  wire[31:0] T48;
  wire[31:0] T49;
  reg [31:0] out_reg_21;
  wire[31:0] T50;
  wire[31:0] T51;
  reg [31:0] out_reg_22;
  wire[31:0] T52;
  wire[31:0] T53;
  reg [31:0] out_reg_23;
  wire[31:0] T54;
  wire[31:0] T55;
  reg [31:0] out_reg_24;
  wire[31:0] T56;
  wire[31:0] T57;
  reg [31:0] out_reg_25;
  wire[31:0] T58;
  wire[31:0] T59;
  reg [31:0] out_reg_26;
  wire[31:0] T60;
  wire[31:0] T61;
  reg [31:0] out_reg_27;
  wire[31:0] T62;
  wire[31:0] T63;
  reg [31:0] out_reg_28;
  wire[31:0] T64;
  wire[31:0] T65;
  reg [31:0] out_reg_29;
  wire[31:0] T66;
  wire[31:0] T67;
  reg [31:0] out_reg_30;
  wire[31:0] T68;
  wire[31:0] T69;
  reg [31:0] out_reg_31;
  wire[31:0] T70;
  wire[31:0] T71;
  reg  start_next_stage_reg;
  wire T74;
  wire T72;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    out_reg_0 = {1{$random}};
    timestamp = {1{$random}};
    out_reg_1 = {1{$random}};
    out_reg_2 = {1{$random}};
    out_reg_3 = {1{$random}};
    out_reg_4 = {1{$random}};
    out_reg_5 = {1{$random}};
    out_reg_6 = {1{$random}};
    out_reg_7 = {1{$random}};
    out_reg_8 = {1{$random}};
    out_reg_9 = {1{$random}};
    out_reg_10 = {1{$random}};
    out_reg_11 = {1{$random}};
    out_reg_12 = {1{$random}};
    out_reg_13 = {1{$random}};
    out_reg_14 = {1{$random}};
    out_reg_15 = {1{$random}};
    out_reg_16 = {1{$random}};
    out_reg_17 = {1{$random}};
    out_reg_18 = {1{$random}};
    out_reg_19 = {1{$random}};
    out_reg_20 = {1{$random}};
    out_reg_21 = {1{$random}};
    out_reg_22 = {1{$random}};
    out_reg_23 = {1{$random}};
    out_reg_24 = {1{$random}};
    out_reg_25 = {1{$random}};
    out_reg_26 = {1{$random}};
    out_reg_27 = {1{$random}};
    out_reg_28 = {1{$random}};
    out_reg_29 = {1{$random}};
    out_reg_30 = {1{$random}};
    out_reg_31 = {1{$random}};
    start_next_stage_reg = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_out_0 = out_reg_0;
  assign T0 = T8 ? io_in_28 : T1;
  assign T1 = T2 ? io_in_0 : out_reg_0;
  assign T2 = T7 & T3;
  assign T3 = timestamp == 1'h0;
  assign T73 = reset ? 1'h0 : T4;
  assign T4 = T6 ? T5 : timestamp;
  assign T5 = timestamp + 1'h1;
  assign T6 = io_clk_en & io_start;
  assign T7 = io_start & io_clk_en;
  assign T8 = T7 & T9;
  assign T9 = timestamp == 1'h1;
  assign io_out_1 = out_reg_1;
  assign T10 = T8 ? io_in_29 : T11;
  assign T11 = T2 ? io_in_1 : out_reg_1;
  assign io_out_2 = out_reg_2;
  assign T12 = T8 ? io_in_30 : T13;
  assign T13 = T2 ? io_in_2 : out_reg_2;
  assign io_out_3 = out_reg_3;
  assign T14 = T8 ? io_in_31 : T15;
  assign T15 = T2 ? io_in_3 : out_reg_3;
  assign io_out_4 = out_reg_4;
  assign T16 = T8 ? io_in_0 : T17;
  assign T17 = T2 ? io_in_4 : out_reg_4;
  assign io_out_5 = out_reg_5;
  assign T18 = T8 ? io_in_1 : T19;
  assign T19 = T2 ? io_in_5 : out_reg_5;
  assign io_out_6 = out_reg_6;
  assign T20 = T8 ? io_in_2 : T21;
  assign T21 = T2 ? io_in_6 : out_reg_6;
  assign io_out_7 = out_reg_7;
  assign T22 = T8 ? io_in_3 : T23;
  assign T23 = T2 ? io_in_7 : out_reg_7;
  assign io_out_8 = out_reg_8;
  assign T24 = T8 ? io_in_4 : T25;
  assign T25 = T2 ? io_in_8 : out_reg_8;
  assign io_out_9 = out_reg_9;
  assign T26 = T8 ? io_in_5 : T27;
  assign T27 = T2 ? io_in_9 : out_reg_9;
  assign io_out_10 = out_reg_10;
  assign T28 = T8 ? io_in_6 : T29;
  assign T29 = T2 ? io_in_10 : out_reg_10;
  assign io_out_11 = out_reg_11;
  assign T30 = T8 ? io_in_7 : T31;
  assign T31 = T2 ? io_in_11 : out_reg_11;
  assign io_out_12 = out_reg_12;
  assign T32 = T8 ? io_in_8 : T33;
  assign T33 = T2 ? io_in_12 : out_reg_12;
  assign io_out_13 = out_reg_13;
  assign T34 = T8 ? io_in_9 : T35;
  assign T35 = T2 ? io_in_13 : out_reg_13;
  assign io_out_14 = out_reg_14;
  assign T36 = T8 ? io_in_10 : T37;
  assign T37 = T2 ? io_in_14 : out_reg_14;
  assign io_out_15 = out_reg_15;
  assign T38 = T8 ? io_in_11 : T39;
  assign T39 = T2 ? io_in_15 : out_reg_15;
  assign io_out_16 = out_reg_16;
  assign T40 = T8 ? io_in_12 : T41;
  assign T41 = T2 ? io_in_16 : out_reg_16;
  assign io_out_17 = out_reg_17;
  assign T42 = T8 ? io_in_13 : T43;
  assign T43 = T2 ? io_in_17 : out_reg_17;
  assign io_out_18 = out_reg_18;
  assign T44 = T8 ? io_in_14 : T45;
  assign T45 = T2 ? io_in_18 : out_reg_18;
  assign io_out_19 = out_reg_19;
  assign T46 = T8 ? io_in_15 : T47;
  assign T47 = T2 ? io_in_19 : out_reg_19;
  assign io_out_20 = out_reg_20;
  assign T48 = T8 ? io_in_16 : T49;
  assign T49 = T2 ? io_in_20 : out_reg_20;
  assign io_out_21 = out_reg_21;
  assign T50 = T8 ? io_in_17 : T51;
  assign T51 = T2 ? io_in_21 : out_reg_21;
  assign io_out_22 = out_reg_22;
  assign T52 = T8 ? io_in_18 : T53;
  assign T53 = T2 ? io_in_22 : out_reg_22;
  assign io_out_23 = out_reg_23;
  assign T54 = T8 ? io_in_19 : T55;
  assign T55 = T2 ? io_in_23 : out_reg_23;
  assign io_out_24 = out_reg_24;
  assign T56 = T8 ? io_in_20 : T57;
  assign T57 = T2 ? io_in_24 : out_reg_24;
  assign io_out_25 = out_reg_25;
  assign T58 = T8 ? io_in_21 : T59;
  assign T59 = T2 ? io_in_25 : out_reg_25;
  assign io_out_26 = out_reg_26;
  assign T60 = T8 ? io_in_22 : T61;
  assign T61 = T2 ? io_in_26 : out_reg_26;
  assign io_out_27 = out_reg_27;
  assign T62 = T8 ? io_in_23 : T63;
  assign T63 = T2 ? io_in_27 : out_reg_27;
  assign io_out_28 = out_reg_28;
  assign T64 = T8 ? io_in_24 : T65;
  assign T65 = T2 ? io_in_28 : out_reg_28;
  assign io_out_29 = out_reg_29;
  assign T66 = T8 ? io_in_25 : T67;
  assign T67 = T2 ? io_in_29 : out_reg_29;
  assign io_out_30 = out_reg_30;
  assign T68 = T8 ? io_in_26 : T69;
  assign T69 = T2 ? io_in_30 : out_reg_30;
  assign io_out_31 = out_reg_31;
  assign T70 = T8 ? io_in_27 : T71;
  assign T71 = T2 ? io_in_31 : out_reg_31;
  assign io_start_next_stage = start_next_stage_reg;
  assign T74 = reset ? 1'h0 : T72;
  assign T72 = T6 ? 1'h1 : start_next_stage_reg;

  always @(posedge clk) begin
    if(T8) begin
      out_reg_0 <= io_in_28;
    end else if(T2) begin
      out_reg_0 <= io_in_0;
    end
    if(reset) begin
      timestamp <= 1'h0;
    end else if(T6) begin
      timestamp <= T5;
    end
    if(T8) begin
      out_reg_1 <= io_in_29;
    end else if(T2) begin
      out_reg_1 <= io_in_1;
    end
    if(T8) begin
      out_reg_2 <= io_in_30;
    end else if(T2) begin
      out_reg_2 <= io_in_2;
    end
    if(T8) begin
      out_reg_3 <= io_in_31;
    end else if(T2) begin
      out_reg_3 <= io_in_3;
    end
    if(T8) begin
      out_reg_4 <= io_in_0;
    end else if(T2) begin
      out_reg_4 <= io_in_4;
    end
    if(T8) begin
      out_reg_5 <= io_in_1;
    end else if(T2) begin
      out_reg_5 <= io_in_5;
    end
    if(T8) begin
      out_reg_6 <= io_in_2;
    end else if(T2) begin
      out_reg_6 <= io_in_6;
    end
    if(T8) begin
      out_reg_7 <= io_in_3;
    end else if(T2) begin
      out_reg_7 <= io_in_7;
    end
    if(T8) begin
      out_reg_8 <= io_in_4;
    end else if(T2) begin
      out_reg_8 <= io_in_8;
    end
    if(T8) begin
      out_reg_9 <= io_in_5;
    end else if(T2) begin
      out_reg_9 <= io_in_9;
    end
    if(T8) begin
      out_reg_10 <= io_in_6;
    end else if(T2) begin
      out_reg_10 <= io_in_10;
    end
    if(T8) begin
      out_reg_11 <= io_in_7;
    end else if(T2) begin
      out_reg_11 <= io_in_11;
    end
    if(T8) begin
      out_reg_12 <= io_in_8;
    end else if(T2) begin
      out_reg_12 <= io_in_12;
    end
    if(T8) begin
      out_reg_13 <= io_in_9;
    end else if(T2) begin
      out_reg_13 <= io_in_13;
    end
    if(T8) begin
      out_reg_14 <= io_in_10;
    end else if(T2) begin
      out_reg_14 <= io_in_14;
    end
    if(T8) begin
      out_reg_15 <= io_in_11;
    end else if(T2) begin
      out_reg_15 <= io_in_15;
    end
    if(T8) begin
      out_reg_16 <= io_in_12;
    end else if(T2) begin
      out_reg_16 <= io_in_16;
    end
    if(T8) begin
      out_reg_17 <= io_in_13;
    end else if(T2) begin
      out_reg_17 <= io_in_17;
    end
    if(T8) begin
      out_reg_18 <= io_in_14;
    end else if(T2) begin
      out_reg_18 <= io_in_18;
    end
    if(T8) begin
      out_reg_19 <= io_in_15;
    end else if(T2) begin
      out_reg_19 <= io_in_19;
    end
    if(T8) begin
      out_reg_20 <= io_in_16;
    end else if(T2) begin
      out_reg_20 <= io_in_20;
    end
    if(T8) begin
      out_reg_21 <= io_in_17;
    end else if(T2) begin
      out_reg_21 <= io_in_21;
    end
    if(T8) begin
      out_reg_22 <= io_in_18;
    end else if(T2) begin
      out_reg_22 <= io_in_22;
    end
    if(T8) begin
      out_reg_23 <= io_in_19;
    end else if(T2) begin
      out_reg_23 <= io_in_23;
    end
    if(T8) begin
      out_reg_24 <= io_in_20;
    end else if(T2) begin
      out_reg_24 <= io_in_24;
    end
    if(T8) begin
      out_reg_25 <= io_in_21;
    end else if(T2) begin
      out_reg_25 <= io_in_25;
    end
    if(T8) begin
      out_reg_26 <= io_in_22;
    end else if(T2) begin
      out_reg_26 <= io_in_26;
    end
    if(T8) begin
      out_reg_27 <= io_in_23;
    end else if(T2) begin
      out_reg_27 <= io_in_27;
    end
    if(T8) begin
      out_reg_28 <= io_in_24;
    end else if(T2) begin
      out_reg_28 <= io_in_28;
    end
    if(T8) begin
      out_reg_29 <= io_in_25;
    end else if(T2) begin
      out_reg_29 <= io_in_29;
    end
    if(T8) begin
      out_reg_30 <= io_in_26;
    end else if(T2) begin
      out_reg_30 <= io_in_30;
    end
    if(T8) begin
      out_reg_31 <= io_in_27;
    end else if(T2) begin
      out_reg_31 <= io_in_31;
    end
    if(reset) begin
      start_next_stage_reg <= 1'h0;
    end else if(T6) begin
      start_next_stage_reg <= 1'h1;
    end
  end
endmodule

module single_port_ram(input clk,
    input [31:0] io_data,
    input  io_addr,
    input  io_we,
    output[31:0] io_q
);

  reg [31:0] out;
  wire[31:0] T0;
  wire[31:0] T1;
  reg [31:0] myMem [1:0];
  wire[31:0] T2;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    out = {1{$random}};
    for (initvar = 0; initvar < 2; initvar = initvar+1)
      myMem[initvar] = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_q = out;
  assign T0 = io_we ? T1 : out;
  assign T1 = myMem[io_addr];

  always @(posedge clk) begin
    if(io_we) begin
      out <= T1;
    end
    if (io_we)
      myMem[io_addr] <= io_data;
  end
endmodule

module memArray(input clk, input reset,
    input  io_clk_en,
    input  io_start,
    output io_start_next_stage,
    input [31:0] io_in_31,
    input [31:0] io_in_30,
    input [31:0] io_in_29,
    input [31:0] io_in_28,
    input [31:0] io_in_27,
    input [31:0] io_in_26,
    input [31:0] io_in_25,
    input [31:0] io_in_24,
    input [31:0] io_in_23,
    input [31:0] io_in_22,
    input [31:0] io_in_21,
    input [31:0] io_in_20,
    input [31:0] io_in_19,
    input [31:0] io_in_18,
    input [31:0] io_in_17,
    input [31:0] io_in_16,
    input [31:0] io_in_15,
    input [31:0] io_in_14,
    input [31:0] io_in_13,
    input [31:0] io_in_12,
    input [31:0] io_in_11,
    input [31:0] io_in_10,
    input [31:0] io_in_9,
    input [31:0] io_in_8,
    input [31:0] io_in_7,
    input [31:0] io_in_6,
    input [31:0] io_in_5,
    input [31:0] io_in_4,
    input [31:0] io_in_3,
    input [31:0] io_in_2,
    input [31:0] io_in_1,
    input [31:0] io_in_0,
    output[31:0] io_out_31,
    output[31:0] io_out_30,
    output[31:0] io_out_29,
    output[31:0] io_out_28,
    output[31:0] io_out_27,
    output[31:0] io_out_26,
    output[31:0] io_out_25,
    output[31:0] io_out_24,
    output[31:0] io_out_23,
    output[31:0] io_out_22,
    output[31:0] io_out_21,
    output[31:0] io_out_20,
    output[31:0] io_out_19,
    output[31:0] io_out_18,
    output[31:0] io_out_17,
    output[31:0] io_out_16,
    output[31:0] io_out_15,
    output[31:0] io_out_14,
    output[31:0] io_out_13,
    output[31:0] io_out_12,
    output[31:0] io_out_11,
    output[31:0] io_out_10,
    output[31:0] io_out_9,
    output[31:0] io_out_8,
    output[31:0] io_out_7,
    output[31:0] io_out_6,
    output[31:0] io_out_5,
    output[31:0] io_out_4,
    output[31:0] io_out_3,
    output[31:0] io_out_2,
    output[31:0] io_out_1,
    output[31:0] io_out_0
);

  wire T0;
  reg  address_7;
  wire T121;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  reg [1:0] state;
  wire[1:0] T122;
  wire[1:0] T9;
  wire[1:0] T10;
  wire[1:0] T11;
  wire T12;
  wire T13;
  wire T14;
  reg  counter;
  wire T123;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  reg  address_6;
  wire T124;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  reg  address_5;
  wire T125;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  reg  address_4;
  wire T126;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  reg  address_3;
  wire T127;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  reg  address_2;
  wire T128;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  reg  address_1;
  wire T129;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  reg  address_0;
  wire T130;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  reg  start_next_stage_reg;
  wire T131;
  wire T120;
  wire[31:0] single_port_ram_io_q;
  wire[31:0] single_port_ram_1_io_q;
  wire[31:0] single_port_ram_2_io_q;
  wire[31:0] single_port_ram_3_io_q;
  wire[31:0] single_port_ram_4_io_q;
  wire[31:0] single_port_ram_5_io_q;
  wire[31:0] single_port_ram_6_io_q;
  wire[31:0] single_port_ram_7_io_q;
  wire[31:0] single_port_ram_8_io_q;
  wire[31:0] single_port_ram_9_io_q;
  wire[31:0] single_port_ram_10_io_q;
  wire[31:0] single_port_ram_11_io_q;
  wire[31:0] single_port_ram_12_io_q;
  wire[31:0] single_port_ram_13_io_q;
  wire[31:0] single_port_ram_14_io_q;
  wire[31:0] single_port_ram_15_io_q;
  wire[31:0] single_port_ram_16_io_q;
  wire[31:0] single_port_ram_17_io_q;
  wire[31:0] single_port_ram_18_io_q;
  wire[31:0] single_port_ram_19_io_q;
  wire[31:0] single_port_ram_20_io_q;
  wire[31:0] single_port_ram_21_io_q;
  wire[31:0] single_port_ram_22_io_q;
  wire[31:0] single_port_ram_23_io_q;
  wire[31:0] single_port_ram_24_io_q;
  wire[31:0] single_port_ram_25_io_q;
  wire[31:0] single_port_ram_26_io_q;
  wire[31:0] single_port_ram_27_io_q;
  wire[31:0] single_port_ram_28_io_q;
  wire[31:0] single_port_ram_29_io_q;
  wire[31:0] single_port_ram_30_io_q;
  wire[31:0] single_port_ram_31_io_q;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    address_7 = {1{$random}};
    state = {1{$random}};
    counter = {1{$random}};
    address_6 = {1{$random}};
    address_5 = {1{$random}};
    address_4 = {1{$random}};
    address_3 = {1{$random}};
    address_2 = {1{$random}};
    address_1 = {1{$random}};
    address_0 = {1{$random}};
    start_next_stage_reg = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = io_start & io_clk_en;
  assign T121 = reset ? 1'h0 : T1;
  assign T1 = T31 ? T30 : T2;
  assign T2 = T28 ? 1'h0 : T3;
  assign T3 = T26 ? T25 : T4;
  assign T4 = T13 ? 1'h1 : T5;
  assign T5 = T7 ? T6 : address_7;
  assign T6 = address_7 + 1'h1;
  assign T7 = T12 & T8;
  assign T8 = state == 2'h0;
  assign T122 = reset ? 2'h0 : T9;
  assign T9 = T28 ? 2'h1 : T10;
  assign T10 = T13 ? 2'h2 : T11;
  assign T11 = T7 ? 2'h1 : state;
  assign T12 = io_clk_en & io_start;
  assign T13 = T23 & T14;
  assign T14 = counter == 1'h1;
  assign T123 = reset ? 1'h0 : T15;
  assign T15 = T21 ? T20 : T16;
  assign T16 = T23 ? T19 : T17;
  assign T17 = T7 ? T18 : counter;
  assign T18 = counter + 1'h1;
  assign T19 = counter + 1'h1;
  assign T20 = counter + 1'h1;
  assign T21 = T12 & T22;
  assign T22 = state == 2'h2;
  assign T23 = T12 & T24;
  assign T24 = state == 2'h1;
  assign T25 = address_7 + 1'h1;
  assign T26 = T23 & T27;
  assign T27 = T14 ^ 1'h1;
  assign T28 = T21 & T29;
  assign T29 = counter == 1'h1;
  assign T30 = address_7 - 1'h1;
  assign T31 = T21 & T32;
  assign T32 = T29 ^ 1'h1;
  assign T33 = io_start & io_clk_en;
  assign T34 = io_start & io_clk_en;
  assign T35 = io_start & io_clk_en;
  assign T36 = io_start & io_clk_en;
  assign T124 = reset ? 1'h0 : T37;
  assign T37 = T31 ? T44 : T38;
  assign T38 = T28 ? 1'h0 : T39;
  assign T39 = T26 ? T43 : T40;
  assign T40 = T13 ? 1'h0 : T41;
  assign T41 = T7 ? T42 : address_6;
  assign T42 = address_6 + 1'h1;
  assign T43 = address_6 + 1'h1;
  assign T44 = address_6 - 1'h1;
  assign T45 = io_start & io_clk_en;
  assign T46 = io_start & io_clk_en;
  assign T47 = io_start & io_clk_en;
  assign T48 = io_start & io_clk_en;
  assign T125 = reset ? 1'h0 : T49;
  assign T49 = T31 ? T56 : T50;
  assign T50 = T28 ? 1'h0 : T51;
  assign T51 = T26 ? T55 : T52;
  assign T52 = T13 ? 1'h1 : T53;
  assign T53 = T7 ? T54 : address_5;
  assign T54 = address_5 + 1'h1;
  assign T55 = address_5 + 1'h1;
  assign T56 = address_5 - 1'h1;
  assign T57 = io_start & io_clk_en;
  assign T58 = io_start & io_clk_en;
  assign T59 = io_start & io_clk_en;
  assign T60 = io_start & io_clk_en;
  assign T126 = reset ? 1'h0 : T61;
  assign T61 = T31 ? T68 : T62;
  assign T62 = T28 ? 1'h0 : T63;
  assign T63 = T26 ? T67 : T64;
  assign T64 = T13 ? 1'h0 : T65;
  assign T65 = T7 ? T66 : address_4;
  assign T66 = address_4 + 1'h1;
  assign T67 = address_4 + 1'h1;
  assign T68 = address_4 - 1'h1;
  assign T69 = io_start & io_clk_en;
  assign T70 = io_start & io_clk_en;
  assign T71 = io_start & io_clk_en;
  assign T72 = io_start & io_clk_en;
  assign T127 = reset ? 1'h0 : T73;
  assign T73 = T31 ? T80 : T74;
  assign T74 = T28 ? 1'h0 : T75;
  assign T75 = T26 ? T79 : T76;
  assign T76 = T13 ? 1'h1 : T77;
  assign T77 = T7 ? T78 : address_3;
  assign T78 = address_3 + 1'h1;
  assign T79 = address_3 + 1'h1;
  assign T80 = address_3 - 1'h1;
  assign T81 = io_start & io_clk_en;
  assign T82 = io_start & io_clk_en;
  assign T83 = io_start & io_clk_en;
  assign T84 = io_start & io_clk_en;
  assign T128 = reset ? 1'h0 : T85;
  assign T85 = T31 ? T92 : T86;
  assign T86 = T28 ? 1'h0 : T87;
  assign T87 = T26 ? T91 : T88;
  assign T88 = T13 ? 1'h0 : T89;
  assign T89 = T7 ? T90 : address_2;
  assign T90 = address_2 + 1'h1;
  assign T91 = address_2 + 1'h1;
  assign T92 = address_2 - 1'h1;
  assign T93 = io_start & io_clk_en;
  assign T94 = io_start & io_clk_en;
  assign T95 = io_start & io_clk_en;
  assign T96 = io_start & io_clk_en;
  assign T129 = reset ? 1'h0 : T97;
  assign T97 = T31 ? T104 : T98;
  assign T98 = T28 ? 1'h0 : T99;
  assign T99 = T26 ? T103 : T100;
  assign T100 = T13 ? 1'h1 : T101;
  assign T101 = T7 ? T102 : address_1;
  assign T102 = address_1 + 1'h1;
  assign T103 = address_1 + 1'h1;
  assign T104 = address_1 - 1'h1;
  assign T105 = io_start & io_clk_en;
  assign T106 = io_start & io_clk_en;
  assign T107 = io_start & io_clk_en;
  assign T108 = io_start & io_clk_en;
  assign T130 = reset ? 1'h0 : T109;
  assign T109 = T31 ? T116 : T110;
  assign T110 = T28 ? 1'h0 : T111;
  assign T111 = T26 ? T115 : T112;
  assign T112 = T13 ? 1'h0 : T113;
  assign T113 = T7 ? T114 : address_0;
  assign T114 = address_0 + 1'h1;
  assign T115 = address_0 + 1'h1;
  assign T116 = address_0 - 1'h1;
  assign T117 = io_start & io_clk_en;
  assign T118 = io_start & io_clk_en;
  assign T119 = io_start & io_clk_en;
  assign io_out_0 = single_port_ram_io_q;
  assign io_out_1 = single_port_ram_1_io_q;
  assign io_out_2 = single_port_ram_2_io_q;
  assign io_out_3 = single_port_ram_3_io_q;
  assign io_out_4 = single_port_ram_4_io_q;
  assign io_out_5 = single_port_ram_5_io_q;
  assign io_out_6 = single_port_ram_6_io_q;
  assign io_out_7 = single_port_ram_7_io_q;
  assign io_out_8 = single_port_ram_8_io_q;
  assign io_out_9 = single_port_ram_9_io_q;
  assign io_out_10 = single_port_ram_10_io_q;
  assign io_out_11 = single_port_ram_11_io_q;
  assign io_out_12 = single_port_ram_12_io_q;
  assign io_out_13 = single_port_ram_13_io_q;
  assign io_out_14 = single_port_ram_14_io_q;
  assign io_out_15 = single_port_ram_15_io_q;
  assign io_out_16 = single_port_ram_16_io_q;
  assign io_out_17 = single_port_ram_17_io_q;
  assign io_out_18 = single_port_ram_18_io_q;
  assign io_out_19 = single_port_ram_19_io_q;
  assign io_out_20 = single_port_ram_20_io_q;
  assign io_out_21 = single_port_ram_21_io_q;
  assign io_out_22 = single_port_ram_22_io_q;
  assign io_out_23 = single_port_ram_23_io_q;
  assign io_out_24 = single_port_ram_24_io_q;
  assign io_out_25 = single_port_ram_25_io_q;
  assign io_out_26 = single_port_ram_26_io_q;
  assign io_out_27 = single_port_ram_27_io_q;
  assign io_out_28 = single_port_ram_28_io_q;
  assign io_out_29 = single_port_ram_29_io_q;
  assign io_out_30 = single_port_ram_30_io_q;
  assign io_out_31 = single_port_ram_31_io_q;
  assign io_start_next_stage = start_next_stage_reg;
  assign T131 = reset ? 1'h0 : T120;
  assign T120 = T21 ? 1'h1 : start_next_stage_reg;
  single_port_ram single_port_ram(.clk(clk),
       .io_data( io_in_0 ),
       .io_addr( address_0 ),
       .io_we( T119 ),
       .io_q( single_port_ram_io_q )
  );
  single_port_ram single_port_ram_1(.clk(clk),
       .io_data( io_in_1 ),
       .io_addr( address_0 ),
       .io_we( T118 ),
       .io_q( single_port_ram_1_io_q )
  );
  single_port_ram single_port_ram_2(.clk(clk),
       .io_data( io_in_2 ),
       .io_addr( address_0 ),
       .io_we( T117 ),
       .io_q( single_port_ram_2_io_q )
  );
  single_port_ram single_port_ram_3(.clk(clk),
       .io_data( io_in_3 ),
       .io_addr( address_0 ),
       .io_we( T108 ),
       .io_q( single_port_ram_3_io_q )
  );
  single_port_ram single_port_ram_4(.clk(clk),
       .io_data( io_in_4 ),
       .io_addr( address_1 ),
       .io_we( T107 ),
       .io_q( single_port_ram_4_io_q )
  );
  single_port_ram single_port_ram_5(.clk(clk),
       .io_data( io_in_5 ),
       .io_addr( address_1 ),
       .io_we( T106 ),
       .io_q( single_port_ram_5_io_q )
  );
  single_port_ram single_port_ram_6(.clk(clk),
       .io_data( io_in_6 ),
       .io_addr( address_1 ),
       .io_we( T105 ),
       .io_q( single_port_ram_6_io_q )
  );
  single_port_ram single_port_ram_7(.clk(clk),
       .io_data( io_in_7 ),
       .io_addr( address_1 ),
       .io_we( T96 ),
       .io_q( single_port_ram_7_io_q )
  );
  single_port_ram single_port_ram_8(.clk(clk),
       .io_data( io_in_8 ),
       .io_addr( address_2 ),
       .io_we( T95 ),
       .io_q( single_port_ram_8_io_q )
  );
  single_port_ram single_port_ram_9(.clk(clk),
       .io_data( io_in_9 ),
       .io_addr( address_2 ),
       .io_we( T94 ),
       .io_q( single_port_ram_9_io_q )
  );
  single_port_ram single_port_ram_10(.clk(clk),
       .io_data( io_in_10 ),
       .io_addr( address_2 ),
       .io_we( T93 ),
       .io_q( single_port_ram_10_io_q )
  );
  single_port_ram single_port_ram_11(.clk(clk),
       .io_data( io_in_11 ),
       .io_addr( address_2 ),
       .io_we( T84 ),
       .io_q( single_port_ram_11_io_q )
  );
  single_port_ram single_port_ram_12(.clk(clk),
       .io_data( io_in_12 ),
       .io_addr( address_3 ),
       .io_we( T83 ),
       .io_q( single_port_ram_12_io_q )
  );
  single_port_ram single_port_ram_13(.clk(clk),
       .io_data( io_in_13 ),
       .io_addr( address_3 ),
       .io_we( T82 ),
       .io_q( single_port_ram_13_io_q )
  );
  single_port_ram single_port_ram_14(.clk(clk),
       .io_data( io_in_14 ),
       .io_addr( address_3 ),
       .io_we( T81 ),
       .io_q( single_port_ram_14_io_q )
  );
  single_port_ram single_port_ram_15(.clk(clk),
       .io_data( io_in_15 ),
       .io_addr( address_3 ),
       .io_we( T72 ),
       .io_q( single_port_ram_15_io_q )
  );
  single_port_ram single_port_ram_16(.clk(clk),
       .io_data( io_in_16 ),
       .io_addr( address_4 ),
       .io_we( T71 ),
       .io_q( single_port_ram_16_io_q )
  );
  single_port_ram single_port_ram_17(.clk(clk),
       .io_data( io_in_17 ),
       .io_addr( address_4 ),
       .io_we( T70 ),
       .io_q( single_port_ram_17_io_q )
  );
  single_port_ram single_port_ram_18(.clk(clk),
       .io_data( io_in_18 ),
       .io_addr( address_4 ),
       .io_we( T69 ),
       .io_q( single_port_ram_18_io_q )
  );
  single_port_ram single_port_ram_19(.clk(clk),
       .io_data( io_in_19 ),
       .io_addr( address_4 ),
       .io_we( T60 ),
       .io_q( single_port_ram_19_io_q )
  );
  single_port_ram single_port_ram_20(.clk(clk),
       .io_data( io_in_20 ),
       .io_addr( address_5 ),
       .io_we( T59 ),
       .io_q( single_port_ram_20_io_q )
  );
  single_port_ram single_port_ram_21(.clk(clk),
       .io_data( io_in_21 ),
       .io_addr( address_5 ),
       .io_we( T58 ),
       .io_q( single_port_ram_21_io_q )
  );
  single_port_ram single_port_ram_22(.clk(clk),
       .io_data( io_in_22 ),
       .io_addr( address_5 ),
       .io_we( T57 ),
       .io_q( single_port_ram_22_io_q )
  );
  single_port_ram single_port_ram_23(.clk(clk),
       .io_data( io_in_23 ),
       .io_addr( address_5 ),
       .io_we( T48 ),
       .io_q( single_port_ram_23_io_q )
  );
  single_port_ram single_port_ram_24(.clk(clk),
       .io_data( io_in_24 ),
       .io_addr( address_6 ),
       .io_we( T47 ),
       .io_q( single_port_ram_24_io_q )
  );
  single_port_ram single_port_ram_25(.clk(clk),
       .io_data( io_in_25 ),
       .io_addr( address_6 ),
       .io_we( T46 ),
       .io_q( single_port_ram_25_io_q )
  );
  single_port_ram single_port_ram_26(.clk(clk),
       .io_data( io_in_26 ),
       .io_addr( address_6 ),
       .io_we( T45 ),
       .io_q( single_port_ram_26_io_q )
  );
  single_port_ram single_port_ram_27(.clk(clk),
       .io_data( io_in_27 ),
       .io_addr( address_6 ),
       .io_we( T36 ),
       .io_q( single_port_ram_27_io_q )
  );
  single_port_ram single_port_ram_28(.clk(clk),
       .io_data( io_in_28 ),
       .io_addr( address_7 ),
       .io_we( T35 ),
       .io_q( single_port_ram_28_io_q )
  );
  single_port_ram single_port_ram_29(.clk(clk),
       .io_data( io_in_29 ),
       .io_addr( address_7 ),
       .io_we( T34 ),
       .io_q( single_port_ram_29_io_q )
  );
  single_port_ram single_port_ram_30(.clk(clk),
       .io_data( io_in_30 ),
       .io_addr( address_7 ),
       .io_we( T33 ),
       .io_q( single_port_ram_30_io_q )
  );
  single_port_ram single_port_ram_31(.clk(clk),
       .io_data( io_in_31 ),
       .io_addr( address_7 ),
       .io_we( T0 ),
       .io_q( single_port_ram_31_io_q )
  );

  always @(posedge clk) begin
    if(reset) begin
      address_7 <= 1'h0;
    end else if(T31) begin
      address_7 <= T30;
    end else if(T28) begin
      address_7 <= 1'h0;
    end else if(T26) begin
      address_7 <= T25;
    end else if(T13) begin
      address_7 <= 1'h1;
    end else if(T7) begin
      address_7 <= T6;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(T28) begin
      state <= 2'h1;
    end else if(T13) begin
      state <= 2'h2;
    end else if(T7) begin
      state <= 2'h1;
    end
    if(reset) begin
      counter <= 1'h0;
    end else if(T21) begin
      counter <= T20;
    end else if(T23) begin
      counter <= T19;
    end else if(T7) begin
      counter <= T18;
    end
    if(reset) begin
      address_6 <= 1'h0;
    end else if(T31) begin
      address_6 <= T44;
    end else if(T28) begin
      address_6 <= 1'h0;
    end else if(T26) begin
      address_6 <= T43;
    end else if(T13) begin
      address_6 <= 1'h0;
    end else if(T7) begin
      address_6 <= T42;
    end
    if(reset) begin
      address_5 <= 1'h0;
    end else if(T31) begin
      address_5 <= T56;
    end else if(T28) begin
      address_5 <= 1'h0;
    end else if(T26) begin
      address_5 <= T55;
    end else if(T13) begin
      address_5 <= 1'h1;
    end else if(T7) begin
      address_5 <= T54;
    end
    if(reset) begin
      address_4 <= 1'h0;
    end else if(T31) begin
      address_4 <= T68;
    end else if(T28) begin
      address_4 <= 1'h0;
    end else if(T26) begin
      address_4 <= T67;
    end else if(T13) begin
      address_4 <= 1'h0;
    end else if(T7) begin
      address_4 <= T66;
    end
    if(reset) begin
      address_3 <= 1'h0;
    end else if(T31) begin
      address_3 <= T80;
    end else if(T28) begin
      address_3 <= 1'h0;
    end else if(T26) begin
      address_3 <= T79;
    end else if(T13) begin
      address_3 <= 1'h1;
    end else if(T7) begin
      address_3 <= T78;
    end
    if(reset) begin
      address_2 <= 1'h0;
    end else if(T31) begin
      address_2 <= T92;
    end else if(T28) begin
      address_2 <= 1'h0;
    end else if(T26) begin
      address_2 <= T91;
    end else if(T13) begin
      address_2 <= 1'h0;
    end else if(T7) begin
      address_2 <= T90;
    end
    if(reset) begin
      address_1 <= 1'h0;
    end else if(T31) begin
      address_1 <= T104;
    end else if(T28) begin
      address_1 <= 1'h0;
    end else if(T26) begin
      address_1 <= T103;
    end else if(T13) begin
      address_1 <= 1'h1;
    end else if(T7) begin
      address_1 <= T102;
    end
    if(reset) begin
      address_0 <= 1'h0;
    end else if(T31) begin
      address_0 <= T116;
    end else if(T28) begin
      address_0 <= 1'h0;
    end else if(T26) begin
      address_0 <= T115;
    end else if(T13) begin
      address_0 <= 1'h0;
    end else if(T7) begin
      address_0 <= T114;
    end
    if(reset) begin
      start_next_stage_reg <= 1'h0;
    end else if(T21) begin
      start_next_stage_reg <= 1'h1;
    end
  end
endmodule

module crossbarShiftUp(input clk, input reset,
    input  io_clk_en,
    input  io_start,
    output io_start_next_stage,
    input [31:0] io_in_31,
    input [31:0] io_in_30,
    input [31:0] io_in_29,
    input [31:0] io_in_28,
    input [31:0] io_in_27,
    input [31:0] io_in_26,
    input [31:0] io_in_25,
    input [31:0] io_in_24,
    input [31:0] io_in_23,
    input [31:0] io_in_22,
    input [31:0] io_in_21,
    input [31:0] io_in_20,
    input [31:0] io_in_19,
    input [31:0] io_in_18,
    input [31:0] io_in_17,
    input [31:0] io_in_16,
    input [31:0] io_in_15,
    input [31:0] io_in_14,
    input [31:0] io_in_13,
    input [31:0] io_in_12,
    input [31:0] io_in_11,
    input [31:0] io_in_10,
    input [31:0] io_in_9,
    input [31:0] io_in_8,
    input [31:0] io_in_7,
    input [31:0] io_in_6,
    input [31:0] io_in_5,
    input [31:0] io_in_4,
    input [31:0] io_in_3,
    input [31:0] io_in_2,
    input [31:0] io_in_1,
    input [31:0] io_in_0,
    output[31:0] io_out_31,
    output[31:0] io_out_30,
    output[31:0] io_out_29,
    output[31:0] io_out_28,
    output[31:0] io_out_27,
    output[31:0] io_out_26,
    output[31:0] io_out_25,
    output[31:0] io_out_24,
    output[31:0] io_out_23,
    output[31:0] io_out_22,
    output[31:0] io_out_21,
    output[31:0] io_out_20,
    output[31:0] io_out_19,
    output[31:0] io_out_18,
    output[31:0] io_out_17,
    output[31:0] io_out_16,
    output[31:0] io_out_15,
    output[31:0] io_out_14,
    output[31:0] io_out_13,
    output[31:0] io_out_12,
    output[31:0] io_out_11,
    output[31:0] io_out_10,
    output[31:0] io_out_9,
    output[31:0] io_out_8,
    output[31:0] io_out_7,
    output[31:0] io_out_6,
    output[31:0] io_out_5,
    output[31:0] io_out_4,
    output[31:0] io_out_3,
    output[31:0] io_out_2,
    output[31:0] io_out_1,
    output[31:0] io_out_0
);

  reg [31:0] out_reg_0;
  wire[31:0] T0;
  wire[31:0] T1;
  wire T2;
  wire T3;
  reg  timestamp;
  wire T73;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  reg [31:0] out_reg_1;
  wire[31:0] T10;
  wire[31:0] T11;
  reg [31:0] out_reg_2;
  wire[31:0] T12;
  wire[31:0] T13;
  reg [31:0] out_reg_3;
  wire[31:0] T14;
  wire[31:0] T15;
  reg [31:0] out_reg_4;
  wire[31:0] T16;
  wire[31:0] T17;
  reg [31:0] out_reg_5;
  wire[31:0] T18;
  wire[31:0] T19;
  reg [31:0] out_reg_6;
  wire[31:0] T20;
  wire[31:0] T21;
  reg [31:0] out_reg_7;
  wire[31:0] T22;
  wire[31:0] T23;
  reg [31:0] out_reg_8;
  wire[31:0] T24;
  wire[31:0] T25;
  reg [31:0] out_reg_9;
  wire[31:0] T26;
  wire[31:0] T27;
  reg [31:0] out_reg_10;
  wire[31:0] T28;
  wire[31:0] T29;
  reg [31:0] out_reg_11;
  wire[31:0] T30;
  wire[31:0] T31;
  reg [31:0] out_reg_12;
  wire[31:0] T32;
  wire[31:0] T33;
  reg [31:0] out_reg_13;
  wire[31:0] T34;
  wire[31:0] T35;
  reg [31:0] out_reg_14;
  wire[31:0] T36;
  wire[31:0] T37;
  reg [31:0] out_reg_15;
  wire[31:0] T38;
  wire[31:0] T39;
  reg [31:0] out_reg_16;
  wire[31:0] T40;
  wire[31:0] T41;
  reg [31:0] out_reg_17;
  wire[31:0] T42;
  wire[31:0] T43;
  reg [31:0] out_reg_18;
  wire[31:0] T44;
  wire[31:0] T45;
  reg [31:0] out_reg_19;
  wire[31:0] T46;
  wire[31:0] T47;
  reg [31:0] out_reg_20;
  wire[31:0] T48;
  wire[31:0] T49;
  reg [31:0] out_reg_21;
  wire[31:0] T50;
  wire[31:0] T51;
  reg [31:0] out_reg_22;
  wire[31:0] T52;
  wire[31:0] T53;
  reg [31:0] out_reg_23;
  wire[31:0] T54;
  wire[31:0] T55;
  reg [31:0] out_reg_24;
  wire[31:0] T56;
  wire[31:0] T57;
  reg [31:0] out_reg_25;
  wire[31:0] T58;
  wire[31:0] T59;
  reg [31:0] out_reg_26;
  wire[31:0] T60;
  wire[31:0] T61;
  reg [31:0] out_reg_27;
  wire[31:0] T62;
  wire[31:0] T63;
  reg [31:0] out_reg_28;
  wire[31:0] T64;
  wire[31:0] T65;
  reg [31:0] out_reg_29;
  wire[31:0] T66;
  wire[31:0] T67;
  reg [31:0] out_reg_30;
  wire[31:0] T68;
  wire[31:0] T69;
  reg [31:0] out_reg_31;
  wire[31:0] T70;
  wire[31:0] T71;
  reg  start_next_stage_reg;
  wire T74;
  wire T72;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    out_reg_0 = {1{$random}};
    timestamp = {1{$random}};
    out_reg_1 = {1{$random}};
    out_reg_2 = {1{$random}};
    out_reg_3 = {1{$random}};
    out_reg_4 = {1{$random}};
    out_reg_5 = {1{$random}};
    out_reg_6 = {1{$random}};
    out_reg_7 = {1{$random}};
    out_reg_8 = {1{$random}};
    out_reg_9 = {1{$random}};
    out_reg_10 = {1{$random}};
    out_reg_11 = {1{$random}};
    out_reg_12 = {1{$random}};
    out_reg_13 = {1{$random}};
    out_reg_14 = {1{$random}};
    out_reg_15 = {1{$random}};
    out_reg_16 = {1{$random}};
    out_reg_17 = {1{$random}};
    out_reg_18 = {1{$random}};
    out_reg_19 = {1{$random}};
    out_reg_20 = {1{$random}};
    out_reg_21 = {1{$random}};
    out_reg_22 = {1{$random}};
    out_reg_23 = {1{$random}};
    out_reg_24 = {1{$random}};
    out_reg_25 = {1{$random}};
    out_reg_26 = {1{$random}};
    out_reg_27 = {1{$random}};
    out_reg_28 = {1{$random}};
    out_reg_29 = {1{$random}};
    out_reg_30 = {1{$random}};
    out_reg_31 = {1{$random}};
    start_next_stage_reg = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_out_0 = out_reg_0;
  assign T0 = T8 ? io_in_4 : T1;
  assign T1 = T2 ? io_in_0 : out_reg_0;
  assign T2 = T7 & T3;
  assign T3 = timestamp == 1'h0;
  assign T73 = reset ? 1'h0 : T4;
  assign T4 = T6 ? T5 : timestamp;
  assign T5 = timestamp + 1'h1;
  assign T6 = io_clk_en & io_start;
  assign T7 = io_start & io_clk_en;
  assign T8 = T7 & T9;
  assign T9 = timestamp == 1'h1;
  assign io_out_1 = out_reg_1;
  assign T10 = T8 ? io_in_5 : T11;
  assign T11 = T2 ? io_in_1 : out_reg_1;
  assign io_out_2 = out_reg_2;
  assign T12 = T8 ? io_in_6 : T13;
  assign T13 = T2 ? io_in_2 : out_reg_2;
  assign io_out_3 = out_reg_3;
  assign T14 = T8 ? io_in_7 : T15;
  assign T15 = T2 ? io_in_3 : out_reg_3;
  assign io_out_4 = out_reg_4;
  assign T16 = T8 ? io_in_8 : T17;
  assign T17 = T2 ? io_in_4 : out_reg_4;
  assign io_out_5 = out_reg_5;
  assign T18 = T8 ? io_in_9 : T19;
  assign T19 = T2 ? io_in_5 : out_reg_5;
  assign io_out_6 = out_reg_6;
  assign T20 = T8 ? io_in_10 : T21;
  assign T21 = T2 ? io_in_6 : out_reg_6;
  assign io_out_7 = out_reg_7;
  assign T22 = T8 ? io_in_11 : T23;
  assign T23 = T2 ? io_in_7 : out_reg_7;
  assign io_out_8 = out_reg_8;
  assign T24 = T8 ? io_in_12 : T25;
  assign T25 = T2 ? io_in_8 : out_reg_8;
  assign io_out_9 = out_reg_9;
  assign T26 = T8 ? io_in_13 : T27;
  assign T27 = T2 ? io_in_9 : out_reg_9;
  assign io_out_10 = out_reg_10;
  assign T28 = T8 ? io_in_14 : T29;
  assign T29 = T2 ? io_in_10 : out_reg_10;
  assign io_out_11 = out_reg_11;
  assign T30 = T8 ? io_in_15 : T31;
  assign T31 = T2 ? io_in_11 : out_reg_11;
  assign io_out_12 = out_reg_12;
  assign T32 = T8 ? io_in_16 : T33;
  assign T33 = T2 ? io_in_12 : out_reg_12;
  assign io_out_13 = out_reg_13;
  assign T34 = T8 ? io_in_17 : T35;
  assign T35 = T2 ? io_in_13 : out_reg_13;
  assign io_out_14 = out_reg_14;
  assign T36 = T8 ? io_in_18 : T37;
  assign T37 = T2 ? io_in_14 : out_reg_14;
  assign io_out_15 = out_reg_15;
  assign T38 = T8 ? io_in_19 : T39;
  assign T39 = T2 ? io_in_15 : out_reg_15;
  assign io_out_16 = out_reg_16;
  assign T40 = T8 ? io_in_20 : T41;
  assign T41 = T2 ? io_in_16 : out_reg_16;
  assign io_out_17 = out_reg_17;
  assign T42 = T8 ? io_in_21 : T43;
  assign T43 = T2 ? io_in_17 : out_reg_17;
  assign io_out_18 = out_reg_18;
  assign T44 = T8 ? io_in_22 : T45;
  assign T45 = T2 ? io_in_18 : out_reg_18;
  assign io_out_19 = out_reg_19;
  assign T46 = T8 ? io_in_23 : T47;
  assign T47 = T2 ? io_in_19 : out_reg_19;
  assign io_out_20 = out_reg_20;
  assign T48 = T8 ? io_in_24 : T49;
  assign T49 = T2 ? io_in_20 : out_reg_20;
  assign io_out_21 = out_reg_21;
  assign T50 = T8 ? io_in_25 : T51;
  assign T51 = T2 ? io_in_21 : out_reg_21;
  assign io_out_22 = out_reg_22;
  assign T52 = T8 ? io_in_26 : T53;
  assign T53 = T2 ? io_in_22 : out_reg_22;
  assign io_out_23 = out_reg_23;
  assign T54 = T8 ? io_in_27 : T55;
  assign T55 = T2 ? io_in_23 : out_reg_23;
  assign io_out_24 = out_reg_24;
  assign T56 = T8 ? io_in_28 : T57;
  assign T57 = T2 ? io_in_24 : out_reg_24;
  assign io_out_25 = out_reg_25;
  assign T58 = T8 ? io_in_29 : T59;
  assign T59 = T2 ? io_in_25 : out_reg_25;
  assign io_out_26 = out_reg_26;
  assign T60 = T8 ? io_in_30 : T61;
  assign T61 = T2 ? io_in_26 : out_reg_26;
  assign io_out_27 = out_reg_27;
  assign T62 = T8 ? io_in_31 : T63;
  assign T63 = T2 ? io_in_27 : out_reg_27;
  assign io_out_28 = out_reg_28;
  assign T64 = T8 ? io_in_0 : T65;
  assign T65 = T2 ? io_in_28 : out_reg_28;
  assign io_out_29 = out_reg_29;
  assign T66 = T8 ? io_in_1 : T67;
  assign T67 = T2 ? io_in_29 : out_reg_29;
  assign io_out_30 = out_reg_30;
  assign T68 = T8 ? io_in_2 : T69;
  assign T69 = T2 ? io_in_30 : out_reg_30;
  assign io_out_31 = out_reg_31;
  assign T70 = T8 ? io_in_3 : T71;
  assign T71 = T2 ? io_in_31 : out_reg_31;
  assign io_start_next_stage = start_next_stage_reg;
  assign T74 = reset ? 1'h0 : T72;
  assign T72 = T6 ? 1'h1 : start_next_stage_reg;

  always @(posedge clk) begin
    if(T8) begin
      out_reg_0 <= io_in_4;
    end else if(T2) begin
      out_reg_0 <= io_in_0;
    end
    if(reset) begin
      timestamp <= 1'h0;
    end else if(T6) begin
      timestamp <= T5;
    end
    if(T8) begin
      out_reg_1 <= io_in_5;
    end else if(T2) begin
      out_reg_1 <= io_in_1;
    end
    if(T8) begin
      out_reg_2 <= io_in_6;
    end else if(T2) begin
      out_reg_2 <= io_in_2;
    end
    if(T8) begin
      out_reg_3 <= io_in_7;
    end else if(T2) begin
      out_reg_3 <= io_in_3;
    end
    if(T8) begin
      out_reg_4 <= io_in_8;
    end else if(T2) begin
      out_reg_4 <= io_in_4;
    end
    if(T8) begin
      out_reg_5 <= io_in_9;
    end else if(T2) begin
      out_reg_5 <= io_in_5;
    end
    if(T8) begin
      out_reg_6 <= io_in_10;
    end else if(T2) begin
      out_reg_6 <= io_in_6;
    end
    if(T8) begin
      out_reg_7 <= io_in_11;
    end else if(T2) begin
      out_reg_7 <= io_in_7;
    end
    if(T8) begin
      out_reg_8 <= io_in_12;
    end else if(T2) begin
      out_reg_8 <= io_in_8;
    end
    if(T8) begin
      out_reg_9 <= io_in_13;
    end else if(T2) begin
      out_reg_9 <= io_in_9;
    end
    if(T8) begin
      out_reg_10 <= io_in_14;
    end else if(T2) begin
      out_reg_10 <= io_in_10;
    end
    if(T8) begin
      out_reg_11 <= io_in_15;
    end else if(T2) begin
      out_reg_11 <= io_in_11;
    end
    if(T8) begin
      out_reg_12 <= io_in_16;
    end else if(T2) begin
      out_reg_12 <= io_in_12;
    end
    if(T8) begin
      out_reg_13 <= io_in_17;
    end else if(T2) begin
      out_reg_13 <= io_in_13;
    end
    if(T8) begin
      out_reg_14 <= io_in_18;
    end else if(T2) begin
      out_reg_14 <= io_in_14;
    end
    if(T8) begin
      out_reg_15 <= io_in_19;
    end else if(T2) begin
      out_reg_15 <= io_in_15;
    end
    if(T8) begin
      out_reg_16 <= io_in_20;
    end else if(T2) begin
      out_reg_16 <= io_in_16;
    end
    if(T8) begin
      out_reg_17 <= io_in_21;
    end else if(T2) begin
      out_reg_17 <= io_in_17;
    end
    if(T8) begin
      out_reg_18 <= io_in_22;
    end else if(T2) begin
      out_reg_18 <= io_in_18;
    end
    if(T8) begin
      out_reg_19 <= io_in_23;
    end else if(T2) begin
      out_reg_19 <= io_in_19;
    end
    if(T8) begin
      out_reg_20 <= io_in_24;
    end else if(T2) begin
      out_reg_20 <= io_in_20;
    end
    if(T8) begin
      out_reg_21 <= io_in_25;
    end else if(T2) begin
      out_reg_21 <= io_in_21;
    end
    if(T8) begin
      out_reg_22 <= io_in_26;
    end else if(T2) begin
      out_reg_22 <= io_in_22;
    end
    if(T8) begin
      out_reg_23 <= io_in_27;
    end else if(T2) begin
      out_reg_23 <= io_in_23;
    end
    if(T8) begin
      out_reg_24 <= io_in_28;
    end else if(T2) begin
      out_reg_24 <= io_in_24;
    end
    if(T8) begin
      out_reg_25 <= io_in_29;
    end else if(T2) begin
      out_reg_25 <= io_in_25;
    end
    if(T8) begin
      out_reg_26 <= io_in_30;
    end else if(T2) begin
      out_reg_26 <= io_in_26;
    end
    if(T8) begin
      out_reg_27 <= io_in_31;
    end else if(T2) begin
      out_reg_27 <= io_in_27;
    end
    if(T8) begin
      out_reg_28 <= io_in_0;
    end else if(T2) begin
      out_reg_28 <= io_in_28;
    end
    if(T8) begin
      out_reg_29 <= io_in_1;
    end else if(T2) begin
      out_reg_29 <= io_in_29;
    end
    if(T8) begin
      out_reg_30 <= io_in_2;
    end else if(T2) begin
      out_reg_30 <= io_in_30;
    end
    if(T8) begin
      out_reg_31 <= io_in_3;
    end else if(T2) begin
      out_reg_31 <= io_in_31;
    end
    if(reset) begin
      start_next_stage_reg <= 1'h0;
    end else if(T6) begin
      start_next_stage_reg <= 1'h1;
    end
  end
endmodule

module streamMatrixTransposeTop(input clk, input reset,
    input  io_clk_en,
    input  io_start,
    output io_start_next_stage,
    input [31:0] io_in_31,
    input [31:0] io_in_30,
    input [31:0] io_in_29,
    input [31:0] io_in_28,
    input [31:0] io_in_27,
    input [31:0] io_in_26,
    input [31:0] io_in_25,
    input [31:0] io_in_24,
    input [31:0] io_in_23,
    input [31:0] io_in_22,
    input [31:0] io_in_21,
    input [31:0] io_in_20,
    input [31:0] io_in_19,
    input [31:0] io_in_18,
    input [31:0] io_in_17,
    input [31:0] io_in_16,
    input [31:0] io_in_15,
    input [31:0] io_in_14,
    input [31:0] io_in_13,
    input [31:0] io_in_12,
    input [31:0] io_in_11,
    input [31:0] io_in_10,
    input [31:0] io_in_9,
    input [31:0] io_in_8,
    input [31:0] io_in_7,
    input [31:0] io_in_6,
    input [31:0] io_in_5,
    input [31:0] io_in_4,
    input [31:0] io_in_3,
    input [31:0] io_in_2,
    input [31:0] io_in_1,
    input [31:0] io_in_0,
    output[31:0] io_out_31,
    output[31:0] io_out_30,
    output[31:0] io_out_29,
    output[31:0] io_out_28,
    output[31:0] io_out_27,
    output[31:0] io_out_26,
    output[31:0] io_out_25,
    output[31:0] io_out_24,
    output[31:0] io_out_23,
    output[31:0] io_out_22,
    output[31:0] io_out_21,
    output[31:0] io_out_20,
    output[31:0] io_out_19,
    output[31:0] io_out_18,
    output[31:0] io_out_17,
    output[31:0] io_out_16,
    output[31:0] io_out_15,
    output[31:0] io_out_14,
    output[31:0] io_out_13,
    output[31:0] io_out_12,
    output[31:0] io_out_11,
    output[31:0] io_out_10,
    output[31:0] io_out_9,
    output[31:0] io_out_8,
    output[31:0] io_out_7,
    output[31:0] io_out_6,
    output[31:0] io_out_5,
    output[31:0] io_out_4,
    output[31:0] io_out_3,
    output[31:0] io_out_2,
    output[31:0] io_out_1,
    output[31:0] io_out_0
);

  wire crossbar_io_start_next_stage;
  wire[31:0] crossbar_io_out_31;
  wire[31:0] crossbar_io_out_30;
  wire[31:0] crossbar_io_out_29;
  wire[31:0] crossbar_io_out_28;
  wire[31:0] crossbar_io_out_27;
  wire[31:0] crossbar_io_out_26;
  wire[31:0] crossbar_io_out_25;
  wire[31:0] crossbar_io_out_24;
  wire[31:0] crossbar_io_out_23;
  wire[31:0] crossbar_io_out_22;
  wire[31:0] crossbar_io_out_21;
  wire[31:0] crossbar_io_out_20;
  wire[31:0] crossbar_io_out_19;
  wire[31:0] crossbar_io_out_18;
  wire[31:0] crossbar_io_out_17;
  wire[31:0] crossbar_io_out_16;
  wire[31:0] crossbar_io_out_15;
  wire[31:0] crossbar_io_out_14;
  wire[31:0] crossbar_io_out_13;
  wire[31:0] crossbar_io_out_12;
  wire[31:0] crossbar_io_out_11;
  wire[31:0] crossbar_io_out_10;
  wire[31:0] crossbar_io_out_9;
  wire[31:0] crossbar_io_out_8;
  wire[31:0] crossbar_io_out_7;
  wire[31:0] crossbar_io_out_6;
  wire[31:0] crossbar_io_out_5;
  wire[31:0] crossbar_io_out_4;
  wire[31:0] crossbar_io_out_3;
  wire[31:0] crossbar_io_out_2;
  wire[31:0] crossbar_io_out_1;
  wire[31:0] crossbar_io_out_0;
  wire crossbarShift_io_start_next_stage;
  wire[31:0] crossbarShift_io_out_31;
  wire[31:0] crossbarShift_io_out_30;
  wire[31:0] crossbarShift_io_out_29;
  wire[31:0] crossbarShift_io_out_28;
  wire[31:0] crossbarShift_io_out_27;
  wire[31:0] crossbarShift_io_out_26;
  wire[31:0] crossbarShift_io_out_25;
  wire[31:0] crossbarShift_io_out_24;
  wire[31:0] crossbarShift_io_out_23;
  wire[31:0] crossbarShift_io_out_22;
  wire[31:0] crossbarShift_io_out_21;
  wire[31:0] crossbarShift_io_out_20;
  wire[31:0] crossbarShift_io_out_19;
  wire[31:0] crossbarShift_io_out_18;
  wire[31:0] crossbarShift_io_out_17;
  wire[31:0] crossbarShift_io_out_16;
  wire[31:0] crossbarShift_io_out_15;
  wire[31:0] crossbarShift_io_out_14;
  wire[31:0] crossbarShift_io_out_13;
  wire[31:0] crossbarShift_io_out_12;
  wire[31:0] crossbarShift_io_out_11;
  wire[31:0] crossbarShift_io_out_10;
  wire[31:0] crossbarShift_io_out_9;
  wire[31:0] crossbarShift_io_out_8;
  wire[31:0] crossbarShift_io_out_7;
  wire[31:0] crossbarShift_io_out_6;
  wire[31:0] crossbarShift_io_out_5;
  wire[31:0] crossbarShift_io_out_4;
  wire[31:0] crossbarShift_io_out_3;
  wire[31:0] crossbarShift_io_out_2;
  wire[31:0] crossbarShift_io_out_1;
  wire[31:0] crossbarShift_io_out_0;
  wire crossbarShift_1_io_start_next_stage;
  wire[31:0] crossbarShift_1_io_out_31;
  wire[31:0] crossbarShift_1_io_out_30;
  wire[31:0] crossbarShift_1_io_out_29;
  wire[31:0] crossbarShift_1_io_out_28;
  wire[31:0] crossbarShift_1_io_out_27;
  wire[31:0] crossbarShift_1_io_out_26;
  wire[31:0] crossbarShift_1_io_out_25;
  wire[31:0] crossbarShift_1_io_out_24;
  wire[31:0] crossbarShift_1_io_out_23;
  wire[31:0] crossbarShift_1_io_out_22;
  wire[31:0] crossbarShift_1_io_out_21;
  wire[31:0] crossbarShift_1_io_out_20;
  wire[31:0] crossbarShift_1_io_out_19;
  wire[31:0] crossbarShift_1_io_out_18;
  wire[31:0] crossbarShift_1_io_out_17;
  wire[31:0] crossbarShift_1_io_out_16;
  wire[31:0] crossbarShift_1_io_out_15;
  wire[31:0] crossbarShift_1_io_out_14;
  wire[31:0] crossbarShift_1_io_out_13;
  wire[31:0] crossbarShift_1_io_out_12;
  wire[31:0] crossbarShift_1_io_out_11;
  wire[31:0] crossbarShift_1_io_out_10;
  wire[31:0] crossbarShift_1_io_out_9;
  wire[31:0] crossbarShift_1_io_out_8;
  wire[31:0] crossbarShift_1_io_out_7;
  wire[31:0] crossbarShift_1_io_out_6;
  wire[31:0] crossbarShift_1_io_out_5;
  wire[31:0] crossbarShift_1_io_out_4;
  wire[31:0] crossbarShift_1_io_out_3;
  wire[31:0] crossbarShift_1_io_out_2;
  wire[31:0] crossbarShift_1_io_out_1;
  wire[31:0] crossbarShift_1_io_out_0;
  wire memArray_io_start_next_stage;
  wire[31:0] memArray_io_out_31;
  wire[31:0] memArray_io_out_30;
  wire[31:0] memArray_io_out_29;
  wire[31:0] memArray_io_out_28;
  wire[31:0] memArray_io_out_27;
  wire[31:0] memArray_io_out_26;
  wire[31:0] memArray_io_out_25;
  wire[31:0] memArray_io_out_24;
  wire[31:0] memArray_io_out_23;
  wire[31:0] memArray_io_out_22;
  wire[31:0] memArray_io_out_21;
  wire[31:0] memArray_io_out_20;
  wire[31:0] memArray_io_out_19;
  wire[31:0] memArray_io_out_18;
  wire[31:0] memArray_io_out_17;
  wire[31:0] memArray_io_out_16;
  wire[31:0] memArray_io_out_15;
  wire[31:0] memArray_io_out_14;
  wire[31:0] memArray_io_out_13;
  wire[31:0] memArray_io_out_12;
  wire[31:0] memArray_io_out_11;
  wire[31:0] memArray_io_out_10;
  wire[31:0] memArray_io_out_9;
  wire[31:0] memArray_io_out_8;
  wire[31:0] memArray_io_out_7;
  wire[31:0] memArray_io_out_6;
  wire[31:0] memArray_io_out_5;
  wire[31:0] memArray_io_out_4;
  wire[31:0] memArray_io_out_3;
  wire[31:0] memArray_io_out_2;
  wire[31:0] memArray_io_out_1;
  wire[31:0] memArray_io_out_0;


  assign io_out_0 = crossbarShift_1_io_out_0;
  assign io_out_1 = crossbarShift_1_io_out_1;
  assign io_out_2 = crossbarShift_1_io_out_2;
  assign io_out_3 = crossbarShift_1_io_out_3;
  assign io_out_4 = crossbarShift_1_io_out_4;
  assign io_out_5 = crossbarShift_1_io_out_5;
  assign io_out_6 = crossbarShift_1_io_out_6;
  assign io_out_7 = crossbarShift_1_io_out_7;
  assign io_out_8 = crossbarShift_1_io_out_8;
  assign io_out_9 = crossbarShift_1_io_out_9;
  assign io_out_10 = crossbarShift_1_io_out_10;
  assign io_out_11 = crossbarShift_1_io_out_11;
  assign io_out_12 = crossbarShift_1_io_out_12;
  assign io_out_13 = crossbarShift_1_io_out_13;
  assign io_out_14 = crossbarShift_1_io_out_14;
  assign io_out_15 = crossbarShift_1_io_out_15;
  assign io_out_16 = crossbarShift_1_io_out_16;
  assign io_out_17 = crossbarShift_1_io_out_17;
  assign io_out_18 = crossbarShift_1_io_out_18;
  assign io_out_19 = crossbarShift_1_io_out_19;
  assign io_out_20 = crossbarShift_1_io_out_20;
  assign io_out_21 = crossbarShift_1_io_out_21;
  assign io_out_22 = crossbarShift_1_io_out_22;
  assign io_out_23 = crossbarShift_1_io_out_23;
  assign io_out_24 = crossbarShift_1_io_out_24;
  assign io_out_25 = crossbarShift_1_io_out_25;
  assign io_out_26 = crossbarShift_1_io_out_26;
  assign io_out_27 = crossbarShift_1_io_out_27;
  assign io_out_28 = crossbarShift_1_io_out_28;
  assign io_out_29 = crossbarShift_1_io_out_29;
  assign io_out_30 = crossbarShift_1_io_out_30;
  assign io_out_31 = crossbarShift_1_io_out_31;
  assign io_start_next_stage = crossbarShift_1_io_start_next_stage;
  crossbar crossbar(.clk(clk), .reset(reset),
       .io_clk_en( io_clk_en ),
       .io_start( io_start ),
       .io_start_next_stage( crossbar_io_start_next_stage ),
       .io_in_31( io_in_31 ),
       .io_in_30( io_in_30 ),
       .io_in_29( io_in_29 ),
       .io_in_28( io_in_28 ),
       .io_in_27( io_in_27 ),
       .io_in_26( io_in_26 ),
       .io_in_25( io_in_25 ),
       .io_in_24( io_in_24 ),
       .io_in_23( io_in_23 ),
       .io_in_22( io_in_22 ),
       .io_in_21( io_in_21 ),
       .io_in_20( io_in_20 ),
       .io_in_19( io_in_19 ),
       .io_in_18( io_in_18 ),
       .io_in_17( io_in_17 ),
       .io_in_16( io_in_16 ),
       .io_in_15( io_in_15 ),
       .io_in_14( io_in_14 ),
       .io_in_13( io_in_13 ),
       .io_in_12( io_in_12 ),
       .io_in_11( io_in_11 ),
       .io_in_10( io_in_10 ),
       .io_in_9( io_in_9 ),
       .io_in_8( io_in_8 ),
       .io_in_7( io_in_7 ),
       .io_in_6( io_in_6 ),
       .io_in_5( io_in_5 ),
       .io_in_4( io_in_4 ),
       .io_in_3( io_in_3 ),
       .io_in_2( io_in_2 ),
       .io_in_1( io_in_1 ),
       .io_in_0( io_in_0 ),
       .io_out_31( crossbar_io_out_31 ),
       .io_out_30( crossbar_io_out_30 ),
       .io_out_29( crossbar_io_out_29 ),
       .io_out_28( crossbar_io_out_28 ),
       .io_out_27( crossbar_io_out_27 ),
       .io_out_26( crossbar_io_out_26 ),
       .io_out_25( crossbar_io_out_25 ),
       .io_out_24( crossbar_io_out_24 ),
       .io_out_23( crossbar_io_out_23 ),
       .io_out_22( crossbar_io_out_22 ),
       .io_out_21( crossbar_io_out_21 ),
       .io_out_20( crossbar_io_out_20 ),
       .io_out_19( crossbar_io_out_19 ),
       .io_out_18( crossbar_io_out_18 ),
       .io_out_17( crossbar_io_out_17 ),
       .io_out_16( crossbar_io_out_16 ),
       .io_out_15( crossbar_io_out_15 ),
       .io_out_14( crossbar_io_out_14 ),
       .io_out_13( crossbar_io_out_13 ),
       .io_out_12( crossbar_io_out_12 ),
       .io_out_11( crossbar_io_out_11 ),
       .io_out_10( crossbar_io_out_10 ),
       .io_out_9( crossbar_io_out_9 ),
       .io_out_8( crossbar_io_out_8 ),
       .io_out_7( crossbar_io_out_7 ),
       .io_out_6( crossbar_io_out_6 ),
       .io_out_5( crossbar_io_out_5 ),
       .io_out_4( crossbar_io_out_4 ),
       .io_out_3( crossbar_io_out_3 ),
       .io_out_2( crossbar_io_out_2 ),
       .io_out_1( crossbar_io_out_1 ),
       .io_out_0( crossbar_io_out_0 )
  );
  crossbarShiftDown crossbarShift(.clk(clk), .reset(reset),
       .io_clk_en( io_clk_en ),
       .io_start( crossbar_io_start_next_stage ),
       .io_start_next_stage( crossbarShift_io_start_next_stage ),
       .io_in_31( crossbar_io_out_31 ),
       .io_in_30( crossbar_io_out_30 ),
       .io_in_29( crossbar_io_out_29 ),
       .io_in_28( crossbar_io_out_28 ),
       .io_in_27( crossbar_io_out_27 ),
       .io_in_26( crossbar_io_out_26 ),
       .io_in_25( crossbar_io_out_25 ),
       .io_in_24( crossbar_io_out_24 ),
       .io_in_23( crossbar_io_out_23 ),
       .io_in_22( crossbar_io_out_22 ),
       .io_in_21( crossbar_io_out_21 ),
       .io_in_20( crossbar_io_out_20 ),
       .io_in_19( crossbar_io_out_19 ),
       .io_in_18( crossbar_io_out_18 ),
       .io_in_17( crossbar_io_out_17 ),
       .io_in_16( crossbar_io_out_16 ),
       .io_in_15( crossbar_io_out_15 ),
       .io_in_14( crossbar_io_out_14 ),
       .io_in_13( crossbar_io_out_13 ),
       .io_in_12( crossbar_io_out_12 ),
       .io_in_11( crossbar_io_out_11 ),
       .io_in_10( crossbar_io_out_10 ),
       .io_in_9( crossbar_io_out_9 ),
       .io_in_8( crossbar_io_out_8 ),
       .io_in_7( crossbar_io_out_7 ),
       .io_in_6( crossbar_io_out_6 ),
       .io_in_5( crossbar_io_out_5 ),
       .io_in_4( crossbar_io_out_4 ),
       .io_in_3( crossbar_io_out_3 ),
       .io_in_2( crossbar_io_out_2 ),
       .io_in_1( crossbar_io_out_1 ),
       .io_in_0( crossbar_io_out_0 ),
       .io_out_31( crossbarShift_io_out_31 ),
       .io_out_30( crossbarShift_io_out_30 ),
       .io_out_29( crossbarShift_io_out_29 ),
       .io_out_28( crossbarShift_io_out_28 ),
       .io_out_27( crossbarShift_io_out_27 ),
       .io_out_26( crossbarShift_io_out_26 ),
       .io_out_25( crossbarShift_io_out_25 ),
       .io_out_24( crossbarShift_io_out_24 ),
       .io_out_23( crossbarShift_io_out_23 ),
       .io_out_22( crossbarShift_io_out_22 ),
       .io_out_21( crossbarShift_io_out_21 ),
       .io_out_20( crossbarShift_io_out_20 ),
       .io_out_19( crossbarShift_io_out_19 ),
       .io_out_18( crossbarShift_io_out_18 ),
       .io_out_17( crossbarShift_io_out_17 ),
       .io_out_16( crossbarShift_io_out_16 ),
       .io_out_15( crossbarShift_io_out_15 ),
       .io_out_14( crossbarShift_io_out_14 ),
       .io_out_13( crossbarShift_io_out_13 ),
       .io_out_12( crossbarShift_io_out_12 ),
       .io_out_11( crossbarShift_io_out_11 ),
       .io_out_10( crossbarShift_io_out_10 ),
       .io_out_9( crossbarShift_io_out_9 ),
       .io_out_8( crossbarShift_io_out_8 ),
       .io_out_7( crossbarShift_io_out_7 ),
       .io_out_6( crossbarShift_io_out_6 ),
       .io_out_5( crossbarShift_io_out_5 ),
       .io_out_4( crossbarShift_io_out_4 ),
       .io_out_3( crossbarShift_io_out_3 ),
       .io_out_2( crossbarShift_io_out_2 ),
       .io_out_1( crossbarShift_io_out_1 ),
       .io_out_0( crossbarShift_io_out_0 )
  );
  memArray memArray(.clk(clk), .reset(reset),
       .io_clk_en( io_clk_en ),
       .io_start( crossbarShift_io_start_next_stage ),
       .io_start_next_stage( memArray_io_start_next_stage ),
       .io_in_31( crossbarShift_io_out_31 ),
       .io_in_30( crossbarShift_io_out_30 ),
       .io_in_29( crossbarShift_io_out_29 ),
       .io_in_28( crossbarShift_io_out_28 ),
       .io_in_27( crossbarShift_io_out_27 ),
       .io_in_26( crossbarShift_io_out_26 ),
       .io_in_25( crossbarShift_io_out_25 ),
       .io_in_24( crossbarShift_io_out_24 ),
       .io_in_23( crossbarShift_io_out_23 ),
       .io_in_22( crossbarShift_io_out_22 ),
       .io_in_21( crossbarShift_io_out_21 ),
       .io_in_20( crossbarShift_io_out_20 ),
       .io_in_19( crossbarShift_io_out_19 ),
       .io_in_18( crossbarShift_io_out_18 ),
       .io_in_17( crossbarShift_io_out_17 ),
       .io_in_16( crossbarShift_io_out_16 ),
       .io_in_15( crossbarShift_io_out_15 ),
       .io_in_14( crossbarShift_io_out_14 ),
       .io_in_13( crossbarShift_io_out_13 ),
       .io_in_12( crossbarShift_io_out_12 ),
       .io_in_11( crossbarShift_io_out_11 ),
       .io_in_10( crossbarShift_io_out_10 ),
       .io_in_9( crossbarShift_io_out_9 ),
       .io_in_8( crossbarShift_io_out_8 ),
       .io_in_7( crossbarShift_io_out_7 ),
       .io_in_6( crossbarShift_io_out_6 ),
       .io_in_5( crossbarShift_io_out_5 ),
       .io_in_4( crossbarShift_io_out_4 ),
       .io_in_3( crossbarShift_io_out_3 ),
       .io_in_2( crossbarShift_io_out_2 ),
       .io_in_1( crossbarShift_io_out_1 ),
       .io_in_0( crossbarShift_io_out_0 ),
       .io_out_31( memArray_io_out_31 ),
       .io_out_30( memArray_io_out_30 ),
       .io_out_29( memArray_io_out_29 ),
       .io_out_28( memArray_io_out_28 ),
       .io_out_27( memArray_io_out_27 ),
       .io_out_26( memArray_io_out_26 ),
       .io_out_25( memArray_io_out_25 ),
       .io_out_24( memArray_io_out_24 ),
       .io_out_23( memArray_io_out_23 ),
       .io_out_22( memArray_io_out_22 ),
       .io_out_21( memArray_io_out_21 ),
       .io_out_20( memArray_io_out_20 ),
       .io_out_19( memArray_io_out_19 ),
       .io_out_18( memArray_io_out_18 ),
       .io_out_17( memArray_io_out_17 ),
       .io_out_16( memArray_io_out_16 ),
       .io_out_15( memArray_io_out_15 ),
       .io_out_14( memArray_io_out_14 ),
       .io_out_13( memArray_io_out_13 ),
       .io_out_12( memArray_io_out_12 ),
       .io_out_11( memArray_io_out_11 ),
       .io_out_10( memArray_io_out_10 ),
       .io_out_9( memArray_io_out_9 ),
       .io_out_8( memArray_io_out_8 ),
       .io_out_7( memArray_io_out_7 ),
       .io_out_6( memArray_io_out_6 ),
       .io_out_5( memArray_io_out_5 ),
       .io_out_4( memArray_io_out_4 ),
       .io_out_3( memArray_io_out_3 ),
       .io_out_2( memArray_io_out_2 ),
       .io_out_1( memArray_io_out_1 ),
       .io_out_0( memArray_io_out_0 )
  );
  crossbarShiftUp crossbarShift_1(.clk(clk), .reset(reset),
       .io_clk_en( io_clk_en ),
       .io_start( memArray_io_start_next_stage ),
       .io_start_next_stage( crossbarShift_1_io_start_next_stage ),
       .io_in_31( memArray_io_out_31 ),
       .io_in_30( memArray_io_out_30 ),
       .io_in_29( memArray_io_out_29 ),
       .io_in_28( memArray_io_out_28 ),
       .io_in_27( memArray_io_out_27 ),
       .io_in_26( memArray_io_out_26 ),
       .io_in_25( memArray_io_out_25 ),
       .io_in_24( memArray_io_out_24 ),
       .io_in_23( memArray_io_out_23 ),
       .io_in_22( memArray_io_out_22 ),
       .io_in_21( memArray_io_out_21 ),
       .io_in_20( memArray_io_out_20 ),
       .io_in_19( memArray_io_out_19 ),
       .io_in_18( memArray_io_out_18 ),
       .io_in_17( memArray_io_out_17 ),
       .io_in_16( memArray_io_out_16 ),
       .io_in_15( memArray_io_out_15 ),
       .io_in_14( memArray_io_out_14 ),
       .io_in_13( memArray_io_out_13 ),
       .io_in_12( memArray_io_out_12 ),
       .io_in_11( memArray_io_out_11 ),
       .io_in_10( memArray_io_out_10 ),
       .io_in_9( memArray_io_out_9 ),
       .io_in_8( memArray_io_out_8 ),
       .io_in_7( memArray_io_out_7 ),
       .io_in_6( memArray_io_out_6 ),
       .io_in_5( memArray_io_out_5 ),
       .io_in_4( memArray_io_out_4 ),
       .io_in_3( memArray_io_out_3 ),
       .io_in_2( memArray_io_out_2 ),
       .io_in_1( memArray_io_out_1 ),
       .io_in_0( memArray_io_out_0 ),
       .io_out_31( crossbarShift_1_io_out_31 ),
       .io_out_30( crossbarShift_1_io_out_30 ),
       .io_out_29( crossbarShift_1_io_out_29 ),
       .io_out_28( crossbarShift_1_io_out_28 ),
       .io_out_27( crossbarShift_1_io_out_27 ),
       .io_out_26( crossbarShift_1_io_out_26 ),
       .io_out_25( crossbarShift_1_io_out_25 ),
       .io_out_24( crossbarShift_1_io_out_24 ),
       .io_out_23( crossbarShift_1_io_out_23 ),
       .io_out_22( crossbarShift_1_io_out_22 ),
       .io_out_21( crossbarShift_1_io_out_21 ),
       .io_out_20( crossbarShift_1_io_out_20 ),
       .io_out_19( crossbarShift_1_io_out_19 ),
       .io_out_18( crossbarShift_1_io_out_18 ),
       .io_out_17( crossbarShift_1_io_out_17 ),
       .io_out_16( crossbarShift_1_io_out_16 ),
       .io_out_15( crossbarShift_1_io_out_15 ),
       .io_out_14( crossbarShift_1_io_out_14 ),
       .io_out_13( crossbarShift_1_io_out_13 ),
       .io_out_12( crossbarShift_1_io_out_12 ),
       .io_out_11( crossbarShift_1_io_out_11 ),
       .io_out_10( crossbarShift_1_io_out_10 ),
       .io_out_9( crossbarShift_1_io_out_9 ),
       .io_out_8( crossbarShift_1_io_out_8 ),
       .io_out_7( crossbarShift_1_io_out_7 ),
       .io_out_6( crossbarShift_1_io_out_6 ),
       .io_out_5( crossbarShift_1_io_out_5 ),
       .io_out_4( crossbarShift_1_io_out_4 ),
       .io_out_3( crossbarShift_1_io_out_3 ),
       .io_out_2( crossbarShift_1_io_out_2 ),
       .io_out_1( crossbarShift_1_io_out_1 ),
       .io_out_0( crossbarShift_1_io_out_0 )
  );
endmodule

module multComplex(input clk, input reset,
    input [15:0] io_real1,
    input [15:0] io_img1,
    input [15:0] io_real2,
    input [15:0] io_img2,
    output[15:0] io_realOut,
    output[15:0] io_imgOut
);

  reg [15:0] delayArrayReal1_1;
  reg [15:0] delayArrayReal1_0;
  reg [15:0] delayArrayImg1_1;
  reg [15:0] delayArrayImg1_0;
  reg [15:0] delayArrayReal2_1;
  reg [15:0] delayArrayReal2_0;
  wire[15:0] addsubfxp_q;
  wire[15:0] addsubfxp_1_q;
  wire[15:0] addsubfxp_2_q;
  wire[15:0] addsubfxp_3_q;
  wire[15:0] addsubfxp_4_q;
  wire[15:0] multfix_q_sc;
  wire[15:0] multfix_1_q_sc;
  wire[15:0] multfix_2_q_sc;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    delayArrayReal1_1 = {1{$random}};
    delayArrayReal1_0 = {1{$random}};
    delayArrayImg1_1 = {1{$random}};
    delayArrayImg1_0 = {1{$random}};
    delayArrayReal2_1 = {1{$random}};
    delayArrayReal2_0 = {1{$random}};
  end
// synthesis translate_on
`endif

  assign io_imgOut = addsubfxp_2_q;
  assign io_realOut = addsubfxp_4_q;
  subfxp # (
    .width(16),
    .cycles(2)
  ) addsubfxp(.clk(clk),
       .a( io_real1 ),
       .b( io_img1 ),
       .q( addsubfxp_q )
  );
  subfxp # (
    .width(16),
    .cycles(2)
  ) addsubfxp_1(.clk(clk),
       .a( io_real2 ),
       .b( io_img2 ),
       .q( addsubfxp_1_q )
  );
  subfxp # (
    .width(16),
    .cycles(2)
  ) addsubfxp_2(.clk(clk),
       .a( multfix_q_sc ),
       .b( multfix_2_q_sc ),
       .q( addsubfxp_2_q )
  );
  addfxp # (
    .width(16),
    .cycles(2)
  ) addsubfxp_3(.clk(clk),
       .a( io_real2 ),
       .b( io_img2 ),
       .q( addsubfxp_3_q )
  );
  addfxp # (
    .width(16),
    .cycles(2)
  ) addsubfxp_4(.clk(clk),
       .a( multfix_q_sc ),
       .b( multfix_1_q_sc ),
       .q( addsubfxp_4_q )
  );
  multfix # (
    .WIDTH(16),
    .CYCLES(1)
  ) multfix(.clk(clk), .rst(reset),
       .a( addsubfxp_q ),
       .b( delayArrayReal2_1 ),
       .q_sc( multfix_q_sc )
       //.q_unsc(  )
  );
  multfix # (
    .WIDTH(16),
    .CYCLES(1)
  ) multfix_1(.clk(clk), .rst(reset),
       .a( delayArrayImg1_1 ),
       .b( addsubfxp_1_q ),
       .q_sc( multfix_1_q_sc )
       //.q_unsc(  )
  );
  multfix # (
    .WIDTH(16),
    .CYCLES(1)
  ) multfix_2(.clk(clk), .rst(reset),
       .a( addsubfxp_3_q ),
       .b( delayArrayReal1_1 ),
       .q_sc( multfix_2_q_sc )
       //.q_unsc(  )
  );

  always @(posedge clk) begin
    delayArrayReal1_1 <= delayArrayReal1_0;
    delayArrayReal1_0 <= io_real1;
    delayArrayImg1_1 <= delayArrayImg1_0;
    delayArrayImg1_0 <= io_img1;
    delayArrayReal2_1 <= delayArrayReal2_0;
    delayArrayReal2_0 <= io_real2;
  end
endmodule

module two_d_convolution(input clk, input reset,
    input  io_clk_en,
    input  io_start,
    output io_start_next_stage,
    input [15:0] io_in_31,
    input [15:0] io_in_30,
    input [15:0] io_in_29,
    input [15:0] io_in_28,
    input [15:0] io_in_27,
    input [15:0] io_in_26,
    input [15:0] io_in_25,
    input [15:0] io_in_24,
    input [15:0] io_in_23,
    input [15:0] io_in_22,
    input [15:0] io_in_21,
    input [15:0] io_in_20,
    input [15:0] io_in_19,
    input [15:0] io_in_18,
    input [15:0] io_in_17,
    input [15:0] io_in_16,
    input [15:0] io_in_15,
    input [15:0] io_in_14,
    input [15:0] io_in_13,
    input [15:0] io_in_12,
    input [15:0] io_in_11,
    input [15:0] io_in_10,
    input [15:0] io_in_9,
    input [15:0] io_in_8,
    input [15:0] io_in_7,
    input [15:0] io_in_6,
    input [15:0] io_in_5,
    input [15:0] io_in_4,
    input [15:0] io_in_3,
    input [15:0] io_in_2,
    input [15:0] io_in_1,
    input [15:0] io_in_0,
    output[15:0] io_out_31,
    output[15:0] io_out_30,
    output[15:0] io_out_29,
    output[15:0] io_out_28,
    output[15:0] io_out_27,
    output[15:0] io_out_26,
    output[15:0] io_out_25,
    output[15:0] io_out_24,
    output[15:0] io_out_23,
    output[15:0] io_out_22,
    output[15:0] io_out_21,
    output[15:0] io_out_20,
    output[15:0] io_out_19,
    output[15:0] io_out_18,
    output[15:0] io_out_17,
    output[15:0] io_out_16,
    output[15:0] io_out_15,
    output[15:0] io_out_14,
    output[15:0] io_out_13,
    output[15:0] io_out_12,
    output[15:0] io_out_11,
    output[15:0] io_out_10,
    output[15:0] io_out_9,
    output[15:0] io_out_8,
    output[15:0] io_out_7,
    output[15:0] io_out_6,
    output[15:0] io_out_5,
    output[15:0] io_out_4,
    output[15:0] io_out_3,
    output[15:0] io_out_2,
    output[15:0] io_out_1,
    output[15:0] io_out_0
);

  wire[31:0] T0;
  wire[31:0] T1;
  wire[31:0] T2;
  wire[31:0] T3;
  wire[31:0] T4;
  wire[31:0] T5;
  wire[31:0] T6;
  wire[31:0] T7;
  wire[31:0] T8;
  wire[31:0] T9;
  wire[31:0] T10;
  wire[31:0] T11;
  wire[31:0] T12;
  wire[31:0] T13;
  wire[31:0] T14;
  wire[31:0] T15;
  wire[31:0] T16;
  wire[31:0] T17;
  wire[31:0] T18;
  wire[31:0] T19;
  wire[31:0] T20;
  wire[31:0] T21;
  wire[31:0] T22;
  wire[31:0] T23;
  wire[31:0] T24;
  wire[31:0] T25;
  wire[31:0] T26;
  wire[31:0] T27;
  wire[31:0] T28;
  wire[31:0] T29;
  wire[31:0] T30;
  wire[31:0] T31;
  reg  startSecondMatrix;
  wire[15:0] T32;
  reg [31:0] delaySecond_24;
  wire[15:0] T33;
  wire[15:0] T34;
  reg [31:0] delaySecond_25;
  wire[15:0] T35;
  wire[15:0] T36;
  reg [31:0] delaySecond_26;
  wire[15:0] T37;
  wire[15:0] T38;
  reg [31:0] delaySecond_27;
  wire[15:0] T39;
  wire[15:0] T40;
  reg [31:0] delaySecond_28;
  wire[15:0] T41;
  wire[15:0] T42;
  reg [31:0] delaySecond_29;
  wire[15:0] T43;
  wire[15:0] T44;
  reg [31:0] delaySecond_30;
  wire[15:0] T45;
  wire[15:0] T46;
  reg [31:0] delaySecond_31;
  wire[15:0] T47;
  wire[15:0] T48;
  reg [31:0] delaySecond_16;
  wire[15:0] T49;
  wire[15:0] T50;
  reg [31:0] delaySecond_17;
  wire[15:0] T51;
  wire[15:0] T52;
  reg [31:0] delaySecond_18;
  wire[15:0] T53;
  wire[15:0] T54;
  reg [31:0] delaySecond_19;
  wire[15:0] T55;
  wire[15:0] T56;
  reg [31:0] delaySecond_20;
  wire[15:0] T57;
  wire[15:0] T58;
  reg [31:0] delaySecond_21;
  wire[15:0] T59;
  wire[15:0] T60;
  reg [31:0] delaySecond_22;
  wire[15:0] T61;
  wire[15:0] T62;
  reg [31:0] delaySecond_23;
  wire[15:0] T63;
  wire[15:0] T64;
  reg [31:0] delaySecond_8;
  wire[15:0] T65;
  wire[15:0] T66;
  reg [31:0] delaySecond_9;
  wire[15:0] T67;
  wire[15:0] T68;
  reg [31:0] delaySecond_10;
  wire[15:0] T69;
  wire[15:0] T70;
  reg [31:0] delaySecond_11;
  wire[15:0] T71;
  wire[15:0] T72;
  reg [31:0] delaySecond_12;
  wire[15:0] T73;
  wire[15:0] T74;
  reg [31:0] delaySecond_13;
  wire[15:0] T75;
  wire[15:0] T76;
  reg [31:0] delaySecond_14;
  wire[15:0] T77;
  wire[15:0] T78;
  reg [31:0] delaySecond_15;
  wire[15:0] T79;
  wire[15:0] T80;
  reg [31:0] delaySecond_0;
  wire[15:0] T81;
  wire[15:0] T82;
  reg [31:0] delaySecond_1;
  wire[15:0] T83;
  wire[15:0] T84;
  reg [31:0] delaySecond_2;
  wire[15:0] T85;
  wire[15:0] T86;
  reg [31:0] delaySecond_3;
  wire[15:0] T87;
  wire[15:0] T88;
  reg [31:0] delaySecond_4;
  wire[15:0] T89;
  wire[15:0] T90;
  reg [31:0] delaySecond_5;
  wire[15:0] T91;
  wire[15:0] T92;
  reg [31:0] delaySecond_6;
  wire[15:0] T93;
  wire[15:0] T94;
  reg [31:0] delaySecond_7;
  wire[15:0] T95;
  reg  delayArrayNext_2;
  reg  delayArrayNext_1;
  reg  delayArrayNext_0;
  wire[15:0] T96;
  reg [31:0] delayFirst_24;
  wire[15:0] T97;
  wire[15:0] T98;
  reg [31:0] delayFirst_25;
  wire[15:0] T99;
  wire[15:0] T100;
  reg [31:0] delayFirst_26;
  wire[15:0] T101;
  wire[15:0] T102;
  reg [31:0] delayFirst_27;
  wire[15:0] T103;
  wire[15:0] T104;
  reg [31:0] delayFirst_28;
  wire[15:0] T105;
  wire[15:0] T106;
  reg [31:0] delayFirst_29;
  wire[15:0] T107;
  wire[15:0] T108;
  reg [31:0] delayFirst_30;
  wire[15:0] T109;
  wire[15:0] T110;
  reg [31:0] delayFirst_31;
  wire[15:0] T111;
  wire[15:0] T112;
  reg [31:0] delayFirst_16;
  wire[15:0] T113;
  wire[15:0] T114;
  reg [31:0] delayFirst_17;
  wire[15:0] T115;
  wire[15:0] T116;
  reg [31:0] delayFirst_18;
  wire[15:0] T117;
  wire[15:0] T118;
  reg [31:0] delayFirst_19;
  wire[15:0] T119;
  wire[15:0] T120;
  reg [31:0] delayFirst_20;
  wire[15:0] T121;
  wire[15:0] T122;
  reg [31:0] delayFirst_21;
  wire[15:0] T123;
  wire[15:0] T124;
  reg [31:0] delayFirst_22;
  wire[15:0] T125;
  wire[15:0] T126;
  reg [31:0] delayFirst_23;
  wire[15:0] T127;
  wire[15:0] T128;
  reg [31:0] delayFirst_8;
  wire[15:0] T129;
  wire[15:0] T130;
  reg [31:0] delayFirst_9;
  wire[15:0] T131;
  wire[15:0] T132;
  reg [31:0] delayFirst_10;
  wire[15:0] T133;
  wire[15:0] T134;
  reg [31:0] delayFirst_11;
  wire[15:0] T135;
  wire[15:0] T136;
  reg [31:0] delayFirst_12;
  wire[15:0] T137;
  wire[15:0] T138;
  reg [31:0] delayFirst_13;
  wire[15:0] T139;
  wire[15:0] T140;
  reg [31:0] delayFirst_14;
  wire[15:0] T141;
  wire[15:0] T142;
  reg [31:0] delayFirst_15;
  wire[15:0] T143;
  wire[15:0] T144;
  reg [31:0] delayFirst_0;
  wire[15:0] T145;
  wire[15:0] T146;
  reg [31:0] delayFirst_1;
  wire[15:0] T147;
  wire[15:0] T148;
  reg [31:0] delayFirst_2;
  wire[15:0] T149;
  wire[15:0] T150;
  reg [31:0] delayFirst_3;
  wire[15:0] T151;
  wire[15:0] T152;
  reg [31:0] delayFirst_4;
  wire[15:0] T153;
  wire[15:0] T154;
  reg [31:0] delayFirst_5;
  wire[15:0] T155;
  wire[15:0] T156;
  reg [31:0] delayFirst_6;
  wire[15:0] T157;
  wire[15:0] T158;
  reg [31:0] delayFirst_7;
  wire[15:0] T159;
  wire[31:0] T160;
  wire[31:0] T161;
  wire[31:0] T162;
  wire[31:0] T163;
  wire[31:0] T164;
  wire[31:0] T165;
  wire[31:0] T166;
  wire[31:0] T167;
  wire[31:0] T168;
  wire[31:0] T169;
  wire[31:0] T170;
  wire[31:0] T171;
  wire[31:0] T172;
  wire[31:0] T173;
  wire[31:0] T174;
  wire[31:0] T175;
  wire[31:0] T176;
  wire[31:0] T177;
  wire[31:0] T178;
  wire[31:0] T179;
  wire[31:0] T180;
  wire[31:0] T181;
  wire[31:0] T182;
  wire[31:0] T183;
  wire[31:0] T184;
  wire[31:0] T185;
  wire[31:0] T186;
  wire[31:0] T187;
  wire[31:0] T188;
  wire[31:0] T189;
  wire[31:0] T190;
  wire[31:0] T191;
  reg  startFirstMatrix;
  reg [15:0] delayInput_24;
  reg [15:0] delayInput_25;
  reg [15:0] delayInput_26;
  reg [15:0] delayInput_27;
  reg [15:0] delayInput_28;
  reg [15:0] delayInput_29;
  reg [15:0] delayInput_30;
  reg [15:0] delayInput_31;
  reg [15:0] delayInput_16;
  reg [15:0] delayInput_17;
  reg [15:0] delayInput_18;
  reg [15:0] delayInput_19;
  reg [15:0] delayInput_20;
  reg [15:0] delayInput_21;
  reg [15:0] delayInput_22;
  reg [15:0] delayInput_23;
  reg [15:0] delayInput_8;
  reg [15:0] delayInput_9;
  reg [15:0] delayInput_10;
  reg [15:0] delayInput_11;
  reg [15:0] delayInput_12;
  reg [15:0] delayInput_13;
  reg [15:0] delayInput_14;
  reg [15:0] delayInput_15;
  reg [15:0] delayInput_0;
  reg [15:0] delayInput_1;
  reg [15:0] delayInput_2;
  reg [15:0] delayInput_3;
  reg [15:0] delayInput_4;
  reg [15:0] delayInput_5;
  reg [15:0] delayInput_6;
  reg [15:0] delayInput_7;
  reg  delayStartNextStage;
  wire fft_next_out;
  wire[15:0] fft_Y15;
  wire[15:0] fft_Y14;
  wire[15:0] fft_Y13;
  wire[15:0] fft_Y12;
  wire[15:0] fft_Y11;
  wire[15:0] fft_Y10;
  wire[15:0] fft_Y9;
  wire[15:0] fft_Y8;
  wire[15:0] fft_Y7;
  wire[15:0] fft_Y6;
  wire[15:0] fft_Y5;
  wire[15:0] fft_Y4;
  wire[15:0] fft_Y3;
  wire[15:0] fft_Y2;
  wire[15:0] fft_Y1;
  wire[15:0] fft_Y0;
  wire[15:0] fft_1_Y15;
  wire[15:0] fft_1_Y14;
  wire[15:0] fft_1_Y13;
  wire[15:0] fft_1_Y12;
  wire[15:0] fft_1_Y11;
  wire[15:0] fft_1_Y10;
  wire[15:0] fft_1_Y9;
  wire[15:0] fft_1_Y8;
  wire[15:0] fft_1_Y7;
  wire[15:0] fft_1_Y6;
  wire[15:0] fft_1_Y5;
  wire[15:0] fft_1_Y4;
  wire[15:0] fft_1_Y3;
  wire[15:0] fft_1_Y2;
  wire[15:0] fft_1_Y1;
  wire[15:0] fft_1_Y0;
  wire[15:0] fft_2_Y15;
  wire[15:0] fft_2_Y14;
  wire[15:0] fft_2_Y13;
  wire[15:0] fft_2_Y12;
  wire[15:0] fft_2_Y11;
  wire[15:0] fft_2_Y10;
  wire[15:0] fft_2_Y9;
  wire[15:0] fft_2_Y8;
  wire[15:0] fft_2_Y7;
  wire[15:0] fft_2_Y6;
  wire[15:0] fft_2_Y5;
  wire[15:0] fft_2_Y4;
  wire[15:0] fft_2_Y3;
  wire[15:0] fft_2_Y2;
  wire[15:0] fft_2_Y1;
  wire[15:0] fft_2_Y0;
  wire[15:0] fft_3_Y15;
  wire[15:0] fft_3_Y14;
  wire[15:0] fft_3_Y13;
  wire[15:0] fft_3_Y12;
  wire[15:0] fft_3_Y11;
  wire[15:0] fft_3_Y10;
  wire[15:0] fft_3_Y9;
  wire[15:0] fft_3_Y8;
  wire[15:0] fft_3_Y7;
  wire[15:0] fft_3_Y6;
  wire[15:0] fft_3_Y5;
  wire[15:0] fft_3_Y4;
  wire[15:0] fft_3_Y3;
  wire[15:0] fft_3_Y2;
  wire[15:0] fft_3_Y1;
  wire[15:0] fft_3_Y0;
  wire fft_4_next_out;
  wire[15:0] fft_4_Y15;
  wire[15:0] fft_4_Y14;
  wire[15:0] fft_4_Y13;
  wire[15:0] fft_4_Y12;
  wire[15:0] fft_4_Y11;
  wire[15:0] fft_4_Y10;
  wire[15:0] fft_4_Y9;
  wire[15:0] fft_4_Y8;
  wire[15:0] fft_4_Y7;
  wire[15:0] fft_4_Y6;
  wire[15:0] fft_4_Y5;
  wire[15:0] fft_4_Y4;
  wire[15:0] fft_4_Y3;
  wire[15:0] fft_4_Y2;
  wire[15:0] fft_4_Y1;
  wire[15:0] fft_4_Y0;
  wire[15:0] fft_5_Y15;
  wire[15:0] fft_5_Y14;
  wire[15:0] fft_5_Y13;
  wire[15:0] fft_5_Y12;
  wire[15:0] fft_5_Y11;
  wire[15:0] fft_5_Y10;
  wire[15:0] fft_5_Y9;
  wire[15:0] fft_5_Y8;
  wire[15:0] fft_5_Y7;
  wire[15:0] fft_5_Y6;
  wire[15:0] fft_5_Y5;
  wire[15:0] fft_5_Y4;
  wire[15:0] fft_5_Y3;
  wire[15:0] fft_5_Y2;
  wire[15:0] fft_5_Y1;
  wire[15:0] fft_5_Y0;
  wire[15:0] fft_6_Y15;
  wire[15:0] fft_6_Y14;
  wire[15:0] fft_6_Y13;
  wire[15:0] fft_6_Y12;
  wire[15:0] fft_6_Y11;
  wire[15:0] fft_6_Y10;
  wire[15:0] fft_6_Y9;
  wire[15:0] fft_6_Y8;
  wire[15:0] fft_6_Y7;
  wire[15:0] fft_6_Y6;
  wire[15:0] fft_6_Y5;
  wire[15:0] fft_6_Y4;
  wire[15:0] fft_6_Y3;
  wire[15:0] fft_6_Y2;
  wire[15:0] fft_6_Y1;
  wire[15:0] fft_6_Y0;
  wire[15:0] fft_7_Y15;
  wire[15:0] fft_7_Y14;
  wire[15:0] fft_7_Y13;
  wire[15:0] fft_7_Y12;
  wire[15:0] fft_7_Y11;
  wire[15:0] fft_7_Y10;
  wire[15:0] fft_7_Y9;
  wire[15:0] fft_7_Y8;
  wire[15:0] fft_7_Y7;
  wire[15:0] fft_7_Y6;
  wire[15:0] fft_7_Y5;
  wire[15:0] fft_7_Y4;
  wire[15:0] fft_7_Y3;
  wire[15:0] fft_7_Y2;
  wire[15:0] fft_7_Y1;
  wire[15:0] fft_7_Y0;
  wire fft_8_next_out;
  wire[15:0] fft_8_Y15;
  wire[15:0] fft_8_Y14;
  wire[15:0] fft_8_Y13;
  wire[15:0] fft_8_Y12;
  wire[15:0] fft_8_Y11;
  wire[15:0] fft_8_Y10;
  wire[15:0] fft_8_Y9;
  wire[15:0] fft_8_Y8;
  wire[15:0] fft_8_Y7;
  wire[15:0] fft_8_Y6;
  wire[15:0] fft_8_Y5;
  wire[15:0] fft_8_Y4;
  wire[15:0] fft_8_Y3;
  wire[15:0] fft_8_Y2;
  wire[15:0] fft_8_Y1;
  wire[15:0] fft_8_Y0;
  wire[15:0] fft_9_Y15;
  wire[15:0] fft_9_Y14;
  wire[15:0] fft_9_Y13;
  wire[15:0] fft_9_Y12;
  wire[15:0] fft_9_Y11;
  wire[15:0] fft_9_Y10;
  wire[15:0] fft_9_Y9;
  wire[15:0] fft_9_Y8;
  wire[15:0] fft_9_Y7;
  wire[15:0] fft_9_Y6;
  wire[15:0] fft_9_Y5;
  wire[15:0] fft_9_Y4;
  wire[15:0] fft_9_Y3;
  wire[15:0] fft_9_Y2;
  wire[15:0] fft_9_Y1;
  wire[15:0] fft_9_Y0;
  wire[15:0] fft_10_Y15;
  wire[15:0] fft_10_Y14;
  wire[15:0] fft_10_Y13;
  wire[15:0] fft_10_Y12;
  wire[15:0] fft_10_Y11;
  wire[15:0] fft_10_Y10;
  wire[15:0] fft_10_Y9;
  wire[15:0] fft_10_Y8;
  wire[15:0] fft_10_Y7;
  wire[15:0] fft_10_Y6;
  wire[15:0] fft_10_Y5;
  wire[15:0] fft_10_Y4;
  wire[15:0] fft_10_Y3;
  wire[15:0] fft_10_Y2;
  wire[15:0] fft_10_Y1;
  wire[15:0] fft_10_Y0;
  wire[15:0] fft_11_Y15;
  wire[15:0] fft_11_Y14;
  wire[15:0] fft_11_Y13;
  wire[15:0] fft_11_Y12;
  wire[15:0] fft_11_Y11;
  wire[15:0] fft_11_Y10;
  wire[15:0] fft_11_Y9;
  wire[15:0] fft_11_Y8;
  wire[15:0] fft_11_Y7;
  wire[15:0] fft_11_Y6;
  wire[15:0] fft_11_Y5;
  wire[15:0] fft_11_Y4;
  wire[15:0] fft_11_Y3;
  wire[15:0] fft_11_Y2;
  wire[15:0] fft_11_Y1;
  wire[15:0] fft_11_Y0;
  wire fft_12_next_out;
  wire[15:0] fft_12_Y14;
  wire[15:0] fft_12_Y12;
  wire[15:0] fft_12_Y10;
  wire[15:0] fft_12_Y8;
  wire[15:0] fft_12_Y6;
  wire[15:0] fft_12_Y4;
  wire[15:0] fft_12_Y2;
  wire[15:0] fft_12_Y0;
  wire[15:0] fft_13_Y14;
  wire[15:0] fft_13_Y12;
  wire[15:0] fft_13_Y10;
  wire[15:0] fft_13_Y8;
  wire[15:0] fft_13_Y6;
  wire[15:0] fft_13_Y4;
  wire[15:0] fft_13_Y2;
  wire[15:0] fft_13_Y0;
  wire[15:0] fft_14_Y14;
  wire[15:0] fft_14_Y12;
  wire[15:0] fft_14_Y10;
  wire[15:0] fft_14_Y8;
  wire[15:0] fft_14_Y6;
  wire[15:0] fft_14_Y4;
  wire[15:0] fft_14_Y2;
  wire[15:0] fft_14_Y0;
  wire[15:0] fft_15_Y14;
  wire[15:0] fft_15_Y12;
  wire[15:0] fft_15_Y10;
  wire[15:0] fft_15_Y8;
  wire[15:0] fft_15_Y6;
  wire[15:0] fft_15_Y4;
  wire[15:0] fft_15_Y2;
  wire[15:0] fft_15_Y0;
  wire[15:0] multComplex_io_realOut;
  wire[15:0] multComplex_io_imgOut;
  wire[15:0] multComplex_1_io_realOut;
  wire[15:0] multComplex_1_io_imgOut;
  wire[15:0] multComplex_2_io_realOut;
  wire[15:0] multComplex_2_io_imgOut;
  wire[15:0] multComplex_3_io_realOut;
  wire[15:0] multComplex_3_io_imgOut;
  wire[15:0] multComplex_4_io_realOut;
  wire[15:0] multComplex_4_io_imgOut;
  wire[15:0] multComplex_5_io_realOut;
  wire[15:0] multComplex_5_io_imgOut;
  wire[15:0] multComplex_6_io_realOut;
  wire[15:0] multComplex_6_io_imgOut;
  wire[15:0] multComplex_7_io_realOut;
  wire[15:0] multComplex_7_io_imgOut;
  wire[15:0] multComplex_8_io_realOut;
  wire[15:0] multComplex_8_io_imgOut;
  wire[15:0] multComplex_9_io_realOut;
  wire[15:0] multComplex_9_io_imgOut;
  wire[15:0] multComplex_10_io_realOut;
  wire[15:0] multComplex_10_io_imgOut;
  wire[15:0] multComplex_11_io_realOut;
  wire[15:0] multComplex_11_io_imgOut;
  wire[15:0] multComplex_12_io_realOut;
  wire[15:0] multComplex_12_io_imgOut;
  wire[15:0] multComplex_13_io_realOut;
  wire[15:0] multComplex_13_io_imgOut;
  wire[15:0] multComplex_14_io_realOut;
  wire[15:0] multComplex_14_io_imgOut;
  wire[15:0] multComplex_15_io_realOut;
  wire[15:0] multComplex_15_io_imgOut;
  wire[15:0] multComplex_16_io_realOut;
  wire[15:0] multComplex_16_io_imgOut;
  wire[15:0] multComplex_17_io_realOut;
  wire[15:0] multComplex_17_io_imgOut;
  wire[15:0] multComplex_18_io_realOut;
  wire[15:0] multComplex_18_io_imgOut;
  wire[15:0] multComplex_19_io_realOut;
  wire[15:0] multComplex_19_io_imgOut;
  wire[15:0] multComplex_20_io_realOut;
  wire[15:0] multComplex_20_io_imgOut;
  wire[15:0] multComplex_21_io_realOut;
  wire[15:0] multComplex_21_io_imgOut;
  wire[15:0] multComplex_22_io_realOut;
  wire[15:0] multComplex_22_io_imgOut;
  wire[15:0] multComplex_23_io_realOut;
  wire[15:0] multComplex_23_io_imgOut;
  wire[15:0] multComplex_24_io_realOut;
  wire[15:0] multComplex_24_io_imgOut;
  wire[15:0] multComplex_25_io_realOut;
  wire[15:0] multComplex_25_io_imgOut;
  wire[15:0] multComplex_26_io_realOut;
  wire[15:0] multComplex_26_io_imgOut;
  wire[15:0] multComplex_27_io_realOut;
  wire[15:0] multComplex_27_io_imgOut;
  wire[15:0] multComplex_28_io_realOut;
  wire[15:0] multComplex_28_io_imgOut;
  wire[15:0] multComplex_29_io_realOut;
  wire[15:0] multComplex_29_io_imgOut;
  wire[15:0] multComplex_30_io_realOut;
  wire[15:0] multComplex_30_io_imgOut;
  wire[15:0] multComplex_31_io_realOut;
  wire[15:0] multComplex_31_io_imgOut;
  wire streamMatrixTransposeTop_io_start_next_stage;
  wire[31:0] streamMatrixTransposeTop_io_out_31;
  wire[31:0] streamMatrixTransposeTop_io_out_30;
  wire[31:0] streamMatrixTransposeTop_io_out_29;
  wire[31:0] streamMatrixTransposeTop_io_out_28;
  wire[31:0] streamMatrixTransposeTop_io_out_27;
  wire[31:0] streamMatrixTransposeTop_io_out_26;
  wire[31:0] streamMatrixTransposeTop_io_out_25;
  wire[31:0] streamMatrixTransposeTop_io_out_24;
  wire[31:0] streamMatrixTransposeTop_io_out_23;
  wire[31:0] streamMatrixTransposeTop_io_out_22;
  wire[31:0] streamMatrixTransposeTop_io_out_21;
  wire[31:0] streamMatrixTransposeTop_io_out_20;
  wire[31:0] streamMatrixTransposeTop_io_out_19;
  wire[31:0] streamMatrixTransposeTop_io_out_18;
  wire[31:0] streamMatrixTransposeTop_io_out_17;
  wire[31:0] streamMatrixTransposeTop_io_out_16;
  wire[31:0] streamMatrixTransposeTop_io_out_15;
  wire[31:0] streamMatrixTransposeTop_io_out_14;
  wire[31:0] streamMatrixTransposeTop_io_out_13;
  wire[31:0] streamMatrixTransposeTop_io_out_12;
  wire[31:0] streamMatrixTransposeTop_io_out_11;
  wire[31:0] streamMatrixTransposeTop_io_out_10;
  wire[31:0] streamMatrixTransposeTop_io_out_9;
  wire[31:0] streamMatrixTransposeTop_io_out_8;
  wire[31:0] streamMatrixTransposeTop_io_out_7;
  wire[31:0] streamMatrixTransposeTop_io_out_6;
  wire[31:0] streamMatrixTransposeTop_io_out_5;
  wire[31:0] streamMatrixTransposeTop_io_out_4;
  wire[31:0] streamMatrixTransposeTop_io_out_3;
  wire[31:0] streamMatrixTransposeTop_io_out_2;
  wire[31:0] streamMatrixTransposeTop_io_out_1;
  wire[31:0] streamMatrixTransposeTop_io_out_0;
  wire streamMatrixTransposeTop_1_io_start_next_stage;
  wire[31:0] streamMatrixTransposeTop_1_io_out_31;
  wire[31:0] streamMatrixTransposeTop_1_io_out_30;
  wire[31:0] streamMatrixTransposeTop_1_io_out_29;
  wire[31:0] streamMatrixTransposeTop_1_io_out_28;
  wire[31:0] streamMatrixTransposeTop_1_io_out_27;
  wire[31:0] streamMatrixTransposeTop_1_io_out_26;
  wire[31:0] streamMatrixTransposeTop_1_io_out_25;
  wire[31:0] streamMatrixTransposeTop_1_io_out_24;
  wire[31:0] streamMatrixTransposeTop_1_io_out_23;
  wire[31:0] streamMatrixTransposeTop_1_io_out_22;
  wire[31:0] streamMatrixTransposeTop_1_io_out_21;
  wire[31:0] streamMatrixTransposeTop_1_io_out_20;
  wire[31:0] streamMatrixTransposeTop_1_io_out_19;
  wire[31:0] streamMatrixTransposeTop_1_io_out_18;
  wire[31:0] streamMatrixTransposeTop_1_io_out_17;
  wire[31:0] streamMatrixTransposeTop_1_io_out_16;
  wire[31:0] streamMatrixTransposeTop_1_io_out_15;
  wire[31:0] streamMatrixTransposeTop_1_io_out_14;
  wire[31:0] streamMatrixTransposeTop_1_io_out_13;
  wire[31:0] streamMatrixTransposeTop_1_io_out_12;
  wire[31:0] streamMatrixTransposeTop_1_io_out_11;
  wire[31:0] streamMatrixTransposeTop_1_io_out_10;
  wire[31:0] streamMatrixTransposeTop_1_io_out_9;
  wire[31:0] streamMatrixTransposeTop_1_io_out_8;
  wire[31:0] streamMatrixTransposeTop_1_io_out_7;
  wire[31:0] streamMatrixTransposeTop_1_io_out_6;
  wire[31:0] streamMatrixTransposeTop_1_io_out_5;
  wire[31:0] streamMatrixTransposeTop_1_io_out_4;
  wire[31:0] streamMatrixTransposeTop_1_io_out_3;
  wire[31:0] streamMatrixTransposeTop_1_io_out_2;
  wire[31:0] streamMatrixTransposeTop_1_io_out_1;
  wire[31:0] streamMatrixTransposeTop_1_io_out_0;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    startSecondMatrix = {1{$random}};
    delaySecond_24 = {1{$random}};
    delaySecond_25 = {1{$random}};
    delaySecond_26 = {1{$random}};
    delaySecond_27 = {1{$random}};
    delaySecond_28 = {1{$random}};
    delaySecond_29 = {1{$random}};
    delaySecond_30 = {1{$random}};
    delaySecond_31 = {1{$random}};
    delaySecond_16 = {1{$random}};
    delaySecond_17 = {1{$random}};
    delaySecond_18 = {1{$random}};
    delaySecond_19 = {1{$random}};
    delaySecond_20 = {1{$random}};
    delaySecond_21 = {1{$random}};
    delaySecond_22 = {1{$random}};
    delaySecond_23 = {1{$random}};
    delaySecond_8 = {1{$random}};
    delaySecond_9 = {1{$random}};
    delaySecond_10 = {1{$random}};
    delaySecond_11 = {1{$random}};
    delaySecond_12 = {1{$random}};
    delaySecond_13 = {1{$random}};
    delaySecond_14 = {1{$random}};
    delaySecond_15 = {1{$random}};
    delaySecond_0 = {1{$random}};
    delaySecond_1 = {1{$random}};
    delaySecond_2 = {1{$random}};
    delaySecond_3 = {1{$random}};
    delaySecond_4 = {1{$random}};
    delaySecond_5 = {1{$random}};
    delaySecond_6 = {1{$random}};
    delaySecond_7 = {1{$random}};
    delayArrayNext_2 = {1{$random}};
    delayArrayNext_1 = {1{$random}};
    delayArrayNext_0 = {1{$random}};
    delayFirst_24 = {1{$random}};
    delayFirst_25 = {1{$random}};
    delayFirst_26 = {1{$random}};
    delayFirst_27 = {1{$random}};
    delayFirst_28 = {1{$random}};
    delayFirst_29 = {1{$random}};
    delayFirst_30 = {1{$random}};
    delayFirst_31 = {1{$random}};
    delayFirst_16 = {1{$random}};
    delayFirst_17 = {1{$random}};
    delayFirst_18 = {1{$random}};
    delayFirst_19 = {1{$random}};
    delayFirst_20 = {1{$random}};
    delayFirst_21 = {1{$random}};
    delayFirst_22 = {1{$random}};
    delayFirst_23 = {1{$random}};
    delayFirst_8 = {1{$random}};
    delayFirst_9 = {1{$random}};
    delayFirst_10 = {1{$random}};
    delayFirst_11 = {1{$random}};
    delayFirst_12 = {1{$random}};
    delayFirst_13 = {1{$random}};
    delayFirst_14 = {1{$random}};
    delayFirst_15 = {1{$random}};
    delayFirst_0 = {1{$random}};
    delayFirst_1 = {1{$random}};
    delayFirst_2 = {1{$random}};
    delayFirst_3 = {1{$random}};
    delayFirst_4 = {1{$random}};
    delayFirst_5 = {1{$random}};
    delayFirst_6 = {1{$random}};
    delayFirst_7 = {1{$random}};
    startFirstMatrix = {1{$random}};
    delayInput_24 = {1{$random}};
    delayInput_25 = {1{$random}};
    delayInput_26 = {1{$random}};
    delayInput_27 = {1{$random}};
    delayInput_28 = {1{$random}};
    delayInput_29 = {1{$random}};
    delayInput_30 = {1{$random}};
    delayInput_31 = {1{$random}};
    delayInput_16 = {1{$random}};
    delayInput_17 = {1{$random}};
    delayInput_18 = {1{$random}};
    delayInput_19 = {1{$random}};
    delayInput_20 = {1{$random}};
    delayInput_21 = {1{$random}};
    delayInput_22 = {1{$random}};
    delayInput_23 = {1{$random}};
    delayInput_8 = {1{$random}};
    delayInput_9 = {1{$random}};
    delayInput_10 = {1{$random}};
    delayInput_11 = {1{$random}};
    delayInput_12 = {1{$random}};
    delayInput_13 = {1{$random}};
    delayInput_14 = {1{$random}};
    delayInput_15 = {1{$random}};
    delayInput_0 = {1{$random}};
    delayInput_1 = {1{$random}};
    delayInput_2 = {1{$random}};
    delayInput_3 = {1{$random}};
    delayInput_4 = {1{$random}};
    delayInput_5 = {1{$random}};
    delayInput_6 = {1{$random}};
    delayInput_7 = {1{$random}};
    delayStartNextStage = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = {fft_8_Y1, fft_8_Y0};
  assign T1 = {fft_8_Y3, fft_8_Y2};
  assign T2 = {fft_8_Y5, fft_8_Y4};
  assign T3 = {fft_8_Y7, fft_8_Y6};
  assign T4 = {fft_8_Y9, fft_8_Y8};
  assign T5 = {fft_8_Y11, fft_8_Y10};
  assign T6 = {fft_8_Y13, fft_8_Y12};
  assign T7 = {fft_8_Y15, fft_8_Y14};
  assign T8 = {fft_9_Y1, fft_9_Y0};
  assign T9 = {fft_9_Y3, fft_9_Y2};
  assign T10 = {fft_9_Y5, fft_9_Y4};
  assign T11 = {fft_9_Y7, fft_9_Y6};
  assign T12 = {fft_9_Y9, fft_9_Y8};
  assign T13 = {fft_9_Y11, fft_9_Y10};
  assign T14 = {fft_9_Y13, fft_9_Y12};
  assign T15 = {fft_9_Y15, fft_9_Y14};
  assign T16 = {fft_10_Y1, fft_10_Y0};
  assign T17 = {fft_10_Y3, fft_10_Y2};
  assign T18 = {fft_10_Y5, fft_10_Y4};
  assign T19 = {fft_10_Y7, fft_10_Y6};
  assign T20 = {fft_10_Y9, fft_10_Y8};
  assign T21 = {fft_10_Y11, fft_10_Y10};
  assign T22 = {fft_10_Y13, fft_10_Y12};
  assign T23 = {fft_10_Y15, fft_10_Y14};
  assign T24 = {fft_11_Y1, fft_11_Y0};
  assign T25 = {fft_11_Y3, fft_11_Y2};
  assign T26 = {fft_11_Y5, fft_11_Y4};
  assign T27 = {fft_11_Y7, fft_11_Y6};
  assign T28 = {fft_11_Y9, fft_11_Y8};
  assign T29 = {fft_11_Y11, fft_11_Y10};
  assign T30 = {fft_11_Y13, fft_11_Y12};
  assign T31 = {fft_11_Y15, fft_11_Y14};
  assign T32 = delaySecond_24[15:0];
  assign T33 = delaySecond_24[31:16];
  assign T34 = delaySecond_25[15:0];
  assign T35 = delaySecond_25[31:16];
  assign T36 = delaySecond_26[15:0];
  assign T37 = delaySecond_26[31:16];
  assign T38 = delaySecond_27[15:0];
  assign T39 = delaySecond_27[31:16];
  assign T40 = delaySecond_28[15:0];
  assign T41 = delaySecond_28[31:16];
  assign T42 = delaySecond_29[15:0];
  assign T43 = delaySecond_29[31:16];
  assign T44 = delaySecond_30[15:0];
  assign T45 = delaySecond_30[31:16];
  assign T46 = delaySecond_31[15:0];
  assign T47 = delaySecond_31[31:16];
  assign T48 = delaySecond_16[15:0];
  assign T49 = delaySecond_16[31:16];
  assign T50 = delaySecond_17[15:0];
  assign T51 = delaySecond_17[31:16];
  assign T52 = delaySecond_18[15:0];
  assign T53 = delaySecond_18[31:16];
  assign T54 = delaySecond_19[15:0];
  assign T55 = delaySecond_19[31:16];
  assign T56 = delaySecond_20[15:0];
  assign T57 = delaySecond_20[31:16];
  assign T58 = delaySecond_21[15:0];
  assign T59 = delaySecond_21[31:16];
  assign T60 = delaySecond_22[15:0];
  assign T61 = delaySecond_22[31:16];
  assign T62 = delaySecond_23[15:0];
  assign T63 = delaySecond_23[31:16];
  assign T64 = delaySecond_8[15:0];
  assign T65 = delaySecond_8[31:16];
  assign T66 = delaySecond_9[15:0];
  assign T67 = delaySecond_9[31:16];
  assign T68 = delaySecond_10[15:0];
  assign T69 = delaySecond_10[31:16];
  assign T70 = delaySecond_11[15:0];
  assign T71 = delaySecond_11[31:16];
  assign T72 = delaySecond_12[15:0];
  assign T73 = delaySecond_12[31:16];
  assign T74 = delaySecond_13[15:0];
  assign T75 = delaySecond_13[31:16];
  assign T76 = delaySecond_14[15:0];
  assign T77 = delaySecond_14[31:16];
  assign T78 = delaySecond_15[15:0];
  assign T79 = delaySecond_15[31:16];
  assign T80 = delaySecond_0[15:0];
  assign T81 = delaySecond_0[31:16];
  assign T82 = delaySecond_1[15:0];
  assign T83 = delaySecond_1[31:16];
  assign T84 = delaySecond_2[15:0];
  assign T85 = delaySecond_2[31:16];
  assign T86 = delaySecond_3[15:0];
  assign T87 = delaySecond_3[31:16];
  assign T88 = delaySecond_4[15:0];
  assign T89 = delaySecond_4[31:16];
  assign T90 = delaySecond_5[15:0];
  assign T91 = delaySecond_5[31:16];
  assign T92 = delaySecond_6[15:0];
  assign T93 = delaySecond_6[31:16];
  assign T94 = delaySecond_7[15:0];
  assign T95 = delaySecond_7[31:16];
  assign T96 = delayFirst_24[15:0];
  assign T97 = delayFirst_24[31:16];
  assign T98 = delayFirst_25[15:0];
  assign T99 = delayFirst_25[31:16];
  assign T100 = delayFirst_26[15:0];
  assign T101 = delayFirst_26[31:16];
  assign T102 = delayFirst_27[15:0];
  assign T103 = delayFirst_27[31:16];
  assign T104 = delayFirst_28[15:0];
  assign T105 = delayFirst_28[31:16];
  assign T106 = delayFirst_29[15:0];
  assign T107 = delayFirst_29[31:16];
  assign T108 = delayFirst_30[15:0];
  assign T109 = delayFirst_30[31:16];
  assign T110 = delayFirst_31[15:0];
  assign T111 = delayFirst_31[31:16];
  assign T112 = delayFirst_16[15:0];
  assign T113 = delayFirst_16[31:16];
  assign T114 = delayFirst_17[15:0];
  assign T115 = delayFirst_17[31:16];
  assign T116 = delayFirst_18[15:0];
  assign T117 = delayFirst_18[31:16];
  assign T118 = delayFirst_19[15:0];
  assign T119 = delayFirst_19[31:16];
  assign T120 = delayFirst_20[15:0];
  assign T121 = delayFirst_20[31:16];
  assign T122 = delayFirst_21[15:0];
  assign T123 = delayFirst_21[31:16];
  assign T124 = delayFirst_22[15:0];
  assign T125 = delayFirst_22[31:16];
  assign T126 = delayFirst_23[15:0];
  assign T127 = delayFirst_23[31:16];
  assign T128 = delayFirst_8[15:0];
  assign T129 = delayFirst_8[31:16];
  assign T130 = delayFirst_9[15:0];
  assign T131 = delayFirst_9[31:16];
  assign T132 = delayFirst_10[15:0];
  assign T133 = delayFirst_10[31:16];
  assign T134 = delayFirst_11[15:0];
  assign T135 = delayFirst_11[31:16];
  assign T136 = delayFirst_12[15:0];
  assign T137 = delayFirst_12[31:16];
  assign T138 = delayFirst_13[15:0];
  assign T139 = delayFirst_13[31:16];
  assign T140 = delayFirst_14[15:0];
  assign T141 = delayFirst_14[31:16];
  assign T142 = delayFirst_15[15:0];
  assign T143 = delayFirst_15[31:16];
  assign T144 = delayFirst_0[15:0];
  assign T145 = delayFirst_0[31:16];
  assign T146 = delayFirst_1[15:0];
  assign T147 = delayFirst_1[31:16];
  assign T148 = delayFirst_2[15:0];
  assign T149 = delayFirst_2[31:16];
  assign T150 = delayFirst_3[15:0];
  assign T151 = delayFirst_3[31:16];
  assign T152 = delayFirst_4[15:0];
  assign T153 = delayFirst_4[31:16];
  assign T154 = delayFirst_5[15:0];
  assign T155 = delayFirst_5[31:16];
  assign T156 = delayFirst_6[15:0];
  assign T157 = delayFirst_6[31:16];
  assign T158 = delayFirst_7[15:0];
  assign T159 = delayFirst_7[31:16];
  assign T160 = {fft_Y1, fft_Y0};
  assign T161 = {fft_Y3, fft_Y2};
  assign T162 = {fft_Y5, fft_Y4};
  assign T163 = {fft_Y7, fft_Y6};
  assign T164 = {fft_Y9, fft_Y8};
  assign T165 = {fft_Y11, fft_Y10};
  assign T166 = {fft_Y13, fft_Y12};
  assign T167 = {fft_Y15, fft_Y14};
  assign T168 = {fft_1_Y1, fft_1_Y0};
  assign T169 = {fft_1_Y3, fft_1_Y2};
  assign T170 = {fft_1_Y5, fft_1_Y4};
  assign T171 = {fft_1_Y7, fft_1_Y6};
  assign T172 = {fft_1_Y9, fft_1_Y8};
  assign T173 = {fft_1_Y11, fft_1_Y10};
  assign T174 = {fft_1_Y13, fft_1_Y12};
  assign T175 = {fft_1_Y15, fft_1_Y14};
  assign T176 = {fft_2_Y1, fft_2_Y0};
  assign T177 = {fft_2_Y3, fft_2_Y2};
  assign T178 = {fft_2_Y5, fft_2_Y4};
  assign T179 = {fft_2_Y7, fft_2_Y6};
  assign T180 = {fft_2_Y9, fft_2_Y8};
  assign T181 = {fft_2_Y11, fft_2_Y10};
  assign T182 = {fft_2_Y13, fft_2_Y12};
  assign T183 = {fft_2_Y15, fft_2_Y14};
  assign T184 = {fft_3_Y1, fft_3_Y0};
  assign T185 = {fft_3_Y3, fft_3_Y2};
  assign T186 = {fft_3_Y5, fft_3_Y4};
  assign T187 = {fft_3_Y7, fft_3_Y6};
  assign T188 = {fft_3_Y9, fft_3_Y8};
  assign T189 = {fft_3_Y11, fft_3_Y10};
  assign T190 = {fft_3_Y13, fft_3_Y12};
  assign T191 = {fft_3_Y15, fft_3_Y14};
  assign io_out_0 = fft_12_Y0;
  assign io_out_1 = fft_12_Y2;
  assign io_out_2 = fft_12_Y4;
  assign io_out_3 = fft_12_Y6;
  assign io_out_4 = fft_12_Y8;
  assign io_out_5 = fft_12_Y10;
  assign io_out_6 = fft_12_Y12;
  assign io_out_7 = fft_12_Y14;
  assign io_out_8 = fft_13_Y0;
  assign io_out_9 = fft_13_Y2;
  assign io_out_10 = fft_13_Y4;
  assign io_out_11 = fft_13_Y6;
  assign io_out_12 = fft_13_Y8;
  assign io_out_13 = fft_13_Y10;
  assign io_out_14 = fft_13_Y12;
  assign io_out_15 = fft_13_Y14;
  assign io_out_16 = fft_14_Y0;
  assign io_out_17 = fft_14_Y2;
  assign io_out_18 = fft_14_Y4;
  assign io_out_19 = fft_14_Y6;
  assign io_out_20 = fft_14_Y8;
  assign io_out_21 = fft_14_Y10;
  assign io_out_22 = fft_14_Y12;
  assign io_out_23 = fft_14_Y14;
  assign io_out_24 = fft_15_Y0;
  assign io_out_25 = fft_15_Y2;
  assign io_out_26 = fft_15_Y4;
  assign io_out_27 = fft_15_Y6;
  assign io_out_28 = fft_15_Y8;
  assign io_out_29 = fft_15_Y10;
  assign io_out_30 = fft_15_Y12;
  assign io_out_31 = fft_15_Y14;
  assign io_start_next_stage = delayStartNextStage;
  fft8_8 fft(.clk(clk), .reset(reset),
       .next( io_start ),
       .next_out( fft_next_out ),
       .X15( 16'h0 ),
       .X14( delayInput_7 ),
       .X13( 16'h0 ),
       .X12( delayInput_6 ),
       .X11( 16'h0 ),
       .X10( delayInput_5 ),
       .X9( 16'h0 ),
       .X8( delayInput_4 ),
       .X7( 16'h0 ),
       .X6( delayInput_3 ),
       .X5( 16'h0 ),
       .X4( delayInput_2 ),
       .X3( 16'h0 ),
       .X2( delayInput_1 ),
       .X1( 16'h0 ),
       .X0( delayInput_0 ),
       .Y15( fft_Y15 ),
       .Y14( fft_Y14 ),
       .Y13( fft_Y13 ),
       .Y12( fft_Y12 ),
       .Y11( fft_Y11 ),
       .Y10( fft_Y10 ),
       .Y9( fft_Y9 ),
       .Y8( fft_Y8 ),
       .Y7( fft_Y7 ),
       .Y6( fft_Y6 ),
       .Y5( fft_Y5 ),
       .Y4( fft_Y4 ),
       .Y3( fft_Y3 ),
       .Y2( fft_Y2 ),
       .Y1( fft_Y1 ),
       .Y0( fft_Y0 )
  );
  fft8_8 fft_1(.clk(clk), .reset(reset),
       .next( io_start ),
       //.next_out(  )
       .X15( 16'h0 ),
       .X14( delayInput_15 ),
       .X13( 16'h0 ),
       .X12( delayInput_14 ),
       .X11( 16'h0 ),
       .X10( delayInput_13 ),
       .X9( 16'h0 ),
       .X8( delayInput_12 ),
       .X7( 16'h0 ),
       .X6( delayInput_11 ),
       .X5( 16'h0 ),
       .X4( delayInput_10 ),
       .X3( 16'h0 ),
       .X2( delayInput_9 ),
       .X1( 16'h0 ),
       .X0( delayInput_8 ),
       .Y15( fft_1_Y15 ),
       .Y14( fft_1_Y14 ),
       .Y13( fft_1_Y13 ),
       .Y12( fft_1_Y12 ),
       .Y11( fft_1_Y11 ),
       .Y10( fft_1_Y10 ),
       .Y9( fft_1_Y9 ),
       .Y8( fft_1_Y8 ),
       .Y7( fft_1_Y7 ),
       .Y6( fft_1_Y6 ),
       .Y5( fft_1_Y5 ),
       .Y4( fft_1_Y4 ),
       .Y3( fft_1_Y3 ),
       .Y2( fft_1_Y2 ),
       .Y1( fft_1_Y1 ),
       .Y0( fft_1_Y0 )
  );
  fft8_8 fft_2(.clk(clk), .reset(reset),
       .next( io_start ),
       //.next_out(  )
       .X15( 16'h0 ),
       .X14( delayInput_23 ),
       .X13( 16'h0 ),
       .X12( delayInput_22 ),
       .X11( 16'h0 ),
       .X10( delayInput_21 ),
       .X9( 16'h0 ),
       .X8( delayInput_20 ),
       .X7( 16'h0 ),
       .X6( delayInput_19 ),
       .X5( 16'h0 ),
       .X4( delayInput_18 ),
       .X3( 16'h0 ),
       .X2( delayInput_17 ),
       .X1( 16'h0 ),
       .X0( delayInput_16 ),
       .Y15( fft_2_Y15 ),
       .Y14( fft_2_Y14 ),
       .Y13( fft_2_Y13 ),
       .Y12( fft_2_Y12 ),
       .Y11( fft_2_Y11 ),
       .Y10( fft_2_Y10 ),
       .Y9( fft_2_Y9 ),
       .Y8( fft_2_Y8 ),
       .Y7( fft_2_Y7 ),
       .Y6( fft_2_Y6 ),
       .Y5( fft_2_Y5 ),
       .Y4( fft_2_Y4 ),
       .Y3( fft_2_Y3 ),
       .Y2( fft_2_Y2 ),
       .Y1( fft_2_Y1 ),
       .Y0( fft_2_Y0 )
  );
  fft8_8 fft_3(.clk(clk), .reset(reset),
       .next( io_start ),
       //.next_out(  )
       .X15( 16'h0 ),
       .X14( delayInput_31 ),
       .X13( 16'h0 ),
       .X12( delayInput_30 ),
       .X11( 16'h0 ),
       .X10( delayInput_29 ),
       .X9( 16'h0 ),
       .X8( delayInput_28 ),
       .X7( 16'h0 ),
       .X6( delayInput_27 ),
       .X5( 16'h0 ),
       .X4( delayInput_26 ),
       .X3( 16'h0 ),
       .X2( delayInput_25 ),
       .X1( 16'h0 ),
       .X0( delayInput_24 ),
       .Y15( fft_3_Y15 ),
       .Y14( fft_3_Y14 ),
       .Y13( fft_3_Y13 ),
       .Y12( fft_3_Y12 ),
       .Y11( fft_3_Y11 ),
       .Y10( fft_3_Y10 ),
       .Y9( fft_3_Y9 ),
       .Y8( fft_3_Y8 ),
       .Y7( fft_3_Y7 ),
       .Y6( fft_3_Y6 ),
       .Y5( fft_3_Y5 ),
       .Y4( fft_3_Y4 ),
       .Y3( fft_3_Y3 ),
       .Y2( fft_3_Y2 ),
       .Y1( fft_3_Y1 ),
       .Y0( fft_3_Y0 )
  );
  streamMatrixTransposeTop streamMatrixTransposeTop(.clk(clk), .reset(reset),
       .io_clk_en( 1'h1 ),
       .io_start( startFirstMatrix ),
       .io_start_next_stage( streamMatrixTransposeTop_io_start_next_stage ),
       .io_in_31( T191 ),
       .io_in_30( T190 ),
       .io_in_29( T189 ),
       .io_in_28( T188 ),
       .io_in_27( T187 ),
       .io_in_26( T186 ),
       .io_in_25( T185 ),
       .io_in_24( T184 ),
       .io_in_23( T183 ),
       .io_in_22( T182 ),
       .io_in_21( T181 ),
       .io_in_20( T180 ),
       .io_in_19( T179 ),
       .io_in_18( T178 ),
       .io_in_17( T177 ),
       .io_in_16( T176 ),
       .io_in_15( T175 ),
       .io_in_14( T174 ),
       .io_in_13( T173 ),
       .io_in_12( T172 ),
       .io_in_11( T171 ),
       .io_in_10( T170 ),
       .io_in_9( T169 ),
       .io_in_8( T168 ),
       .io_in_7( T167 ),
       .io_in_6( T166 ),
       .io_in_5( T165 ),
       .io_in_4( T164 ),
       .io_in_3( T163 ),
       .io_in_2( T162 ),
       .io_in_1( T161 ),
       .io_in_0( T160 ),
       .io_out_31( streamMatrixTransposeTop_io_out_31 ),
       .io_out_30( streamMatrixTransposeTop_io_out_30 ),
       .io_out_29( streamMatrixTransposeTop_io_out_29 ),
       .io_out_28( streamMatrixTransposeTop_io_out_28 ),
       .io_out_27( streamMatrixTransposeTop_io_out_27 ),
       .io_out_26( streamMatrixTransposeTop_io_out_26 ),
       .io_out_25( streamMatrixTransposeTop_io_out_25 ),
       .io_out_24( streamMatrixTransposeTop_io_out_24 ),
       .io_out_23( streamMatrixTransposeTop_io_out_23 ),
       .io_out_22( streamMatrixTransposeTop_io_out_22 ),
       .io_out_21( streamMatrixTransposeTop_io_out_21 ),
       .io_out_20( streamMatrixTransposeTop_io_out_20 ),
       .io_out_19( streamMatrixTransposeTop_io_out_19 ),
       .io_out_18( streamMatrixTransposeTop_io_out_18 ),
       .io_out_17( streamMatrixTransposeTop_io_out_17 ),
       .io_out_16( streamMatrixTransposeTop_io_out_16 ),
       .io_out_15( streamMatrixTransposeTop_io_out_15 ),
       .io_out_14( streamMatrixTransposeTop_io_out_14 ),
       .io_out_13( streamMatrixTransposeTop_io_out_13 ),
       .io_out_12( streamMatrixTransposeTop_io_out_12 ),
       .io_out_11( streamMatrixTransposeTop_io_out_11 ),
       .io_out_10( streamMatrixTransposeTop_io_out_10 ),
       .io_out_9( streamMatrixTransposeTop_io_out_9 ),
       .io_out_8( streamMatrixTransposeTop_io_out_8 ),
       .io_out_7( streamMatrixTransposeTop_io_out_7 ),
       .io_out_6( streamMatrixTransposeTop_io_out_6 ),
       .io_out_5( streamMatrixTransposeTop_io_out_5 ),
       .io_out_4( streamMatrixTransposeTop_io_out_4 ),
       .io_out_3( streamMatrixTransposeTop_io_out_3 ),
       .io_out_2( streamMatrixTransposeTop_io_out_2 ),
       .io_out_1( streamMatrixTransposeTop_io_out_1 ),
       .io_out_0( streamMatrixTransposeTop_io_out_0 )
  );
  fft8_8 fft_4(.clk(clk), .reset(reset),
       .next( streamMatrixTransposeTop_io_start_next_stage ),
       .next_out( fft_4_next_out ),
       .X15( T159 ),
       .X14( T158 ),
       .X13( T157 ),
       .X12( T156 ),
       .X11( T155 ),
       .X10( T154 ),
       .X9( T153 ),
       .X8( T152 ),
       .X7( T151 ),
       .X6( T150 ),
       .X5( T149 ),
       .X4( T148 ),
       .X3( T147 ),
       .X2( T146 ),
       .X1( T145 ),
       .X0( T144 ),
       .Y15( fft_4_Y15 ),
       .Y14( fft_4_Y14 ),
       .Y13( fft_4_Y13 ),
       .Y12( fft_4_Y12 ),
       .Y11( fft_4_Y11 ),
       .Y10( fft_4_Y10 ),
       .Y9( fft_4_Y9 ),
       .Y8( fft_4_Y8 ),
       .Y7( fft_4_Y7 ),
       .Y6( fft_4_Y6 ),
       .Y5( fft_4_Y5 ),
       .Y4( fft_4_Y4 ),
       .Y3( fft_4_Y3 ),
       .Y2( fft_4_Y2 ),
       .Y1( fft_4_Y1 ),
       .Y0( fft_4_Y0 )
  );
  fft8_8 fft_5(.clk(clk), .reset(reset),
       .next( streamMatrixTransposeTop_io_start_next_stage ),
       //.next_out(  )
       .X15( T143 ),
       .X14( T142 ),
       .X13( T141 ),
       .X12( T140 ),
       .X11( T139 ),
       .X10( T138 ),
       .X9( T137 ),
       .X8( T136 ),
       .X7( T135 ),
       .X6( T134 ),
       .X5( T133 ),
       .X4( T132 ),
       .X3( T131 ),
       .X2( T130 ),
       .X1( T129 ),
       .X0( T128 ),
       .Y15( fft_5_Y15 ),
       .Y14( fft_5_Y14 ),
       .Y13( fft_5_Y13 ),
       .Y12( fft_5_Y12 ),
       .Y11( fft_5_Y11 ),
       .Y10( fft_5_Y10 ),
       .Y9( fft_5_Y9 ),
       .Y8( fft_5_Y8 ),
       .Y7( fft_5_Y7 ),
       .Y6( fft_5_Y6 ),
       .Y5( fft_5_Y5 ),
       .Y4( fft_5_Y4 ),
       .Y3( fft_5_Y3 ),
       .Y2( fft_5_Y2 ),
       .Y1( fft_5_Y1 ),
       .Y0( fft_5_Y0 )
  );
  fft8_8 fft_6(.clk(clk), .reset(reset),
       .next( streamMatrixTransposeTop_io_start_next_stage ),
       //.next_out(  )
       .X15( T127 ),
       .X14( T126 ),
       .X13( T125 ),
       .X12( T124 ),
       .X11( T123 ),
       .X10( T122 ),
       .X9( T121 ),
       .X8( T120 ),
       .X7( T119 ),
       .X6( T118 ),
       .X5( T117 ),
       .X4( T116 ),
       .X3( T115 ),
       .X2( T114 ),
       .X1( T113 ),
       .X0( T112 ),
       .Y15( fft_6_Y15 ),
       .Y14( fft_6_Y14 ),
       .Y13( fft_6_Y13 ),
       .Y12( fft_6_Y12 ),
       .Y11( fft_6_Y11 ),
       .Y10( fft_6_Y10 ),
       .Y9( fft_6_Y9 ),
       .Y8( fft_6_Y8 ),
       .Y7( fft_6_Y7 ),
       .Y6( fft_6_Y6 ),
       .Y5( fft_6_Y5 ),
       .Y4( fft_6_Y4 ),
       .Y3( fft_6_Y3 ),
       .Y2( fft_6_Y2 ),
       .Y1( fft_6_Y1 ),
       .Y0( fft_6_Y0 )
  );
  fft8_8 fft_7(.clk(clk), .reset(reset),
       .next( streamMatrixTransposeTop_io_start_next_stage ),
       //.next_out(  )
       .X15( T111 ),
       .X14( T110 ),
       .X13( T109 ),
       .X12( T108 ),
       .X11( T107 ),
       .X10( T106 ),
       .X9( T105 ),
       .X8( T104 ),
       .X7( T103 ),
       .X6( T102 ),
       .X5( T101 ),
       .X4( T100 ),
       .X3( T99 ),
       .X2( T98 ),
       .X1( T97 ),
       .X0( T96 ),
       .Y15( fft_7_Y15 ),
       .Y14( fft_7_Y14 ),
       .Y13( fft_7_Y13 ),
       .Y12( fft_7_Y12 ),
       .Y11( fft_7_Y11 ),
       .Y10( fft_7_Y10 ),
       .Y9( fft_7_Y9 ),
       .Y8( fft_7_Y8 ),
       .Y7( fft_7_Y7 ),
       .Y6( fft_7_Y6 ),
       .Y5( fft_7_Y5 ),
       .Y4( fft_7_Y4 ),
       .Y3( fft_7_Y3 ),
       .Y2( fft_7_Y2 ),
       .Y1( fft_7_Y1 ),
       .Y0( fft_7_Y0 )
  );
  multComplex multComplex(.clk(clk), .reset(reset),
       .io_real1( fft_4_Y0 ),
       .io_img1( fft_4_Y1 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_io_realOut ),
       .io_imgOut( multComplex_io_imgOut )
  );
  multComplex multComplex_1(.clk(clk), .reset(reset),
       .io_real1( fft_4_Y2 ),
       .io_img1( fft_4_Y3 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_1_io_realOut ),
       .io_imgOut( multComplex_1_io_imgOut )
  );
  multComplex multComplex_2(.clk(clk), .reset(reset),
       .io_real1( fft_4_Y4 ),
       .io_img1( fft_4_Y5 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_2_io_realOut ),
       .io_imgOut( multComplex_2_io_imgOut )
  );
  multComplex multComplex_3(.clk(clk), .reset(reset),
       .io_real1( fft_4_Y6 ),
       .io_img1( fft_4_Y7 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_3_io_realOut ),
       .io_imgOut( multComplex_3_io_imgOut )
  );
  multComplex multComplex_4(.clk(clk), .reset(reset),
       .io_real1( fft_4_Y8 ),
       .io_img1( fft_4_Y9 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_4_io_realOut ),
       .io_imgOut( multComplex_4_io_imgOut )
  );
  multComplex multComplex_5(.clk(clk), .reset(reset),
       .io_real1( fft_4_Y10 ),
       .io_img1( fft_4_Y11 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_5_io_realOut ),
       .io_imgOut( multComplex_5_io_imgOut )
  );
  multComplex multComplex_6(.clk(clk), .reset(reset),
       .io_real1( fft_4_Y12 ),
       .io_img1( fft_4_Y13 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_6_io_realOut ),
       .io_imgOut( multComplex_6_io_imgOut )
  );
  multComplex multComplex_7(.clk(clk), .reset(reset),
       .io_real1( fft_4_Y14 ),
       .io_img1( fft_4_Y15 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_7_io_realOut ),
       .io_imgOut( multComplex_7_io_imgOut )
  );
  multComplex multComplex_8(.clk(clk), .reset(reset),
       .io_real1( fft_5_Y0 ),
       .io_img1( fft_5_Y1 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_8_io_realOut ),
       .io_imgOut( multComplex_8_io_imgOut )
  );
  multComplex multComplex_9(.clk(clk), .reset(reset),
       .io_real1( fft_5_Y2 ),
       .io_img1( fft_5_Y3 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_9_io_realOut ),
       .io_imgOut( multComplex_9_io_imgOut )
  );
  multComplex multComplex_10(.clk(clk), .reset(reset),
       .io_real1( fft_5_Y4 ),
       .io_img1( fft_5_Y5 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_10_io_realOut ),
       .io_imgOut( multComplex_10_io_imgOut )
  );
  multComplex multComplex_11(.clk(clk), .reset(reset),
       .io_real1( fft_5_Y6 ),
       .io_img1( fft_5_Y7 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_11_io_realOut ),
       .io_imgOut( multComplex_11_io_imgOut )
  );
  multComplex multComplex_12(.clk(clk), .reset(reset),
       .io_real1( fft_5_Y8 ),
       .io_img1( fft_5_Y9 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_12_io_realOut ),
       .io_imgOut( multComplex_12_io_imgOut )
  );
  multComplex multComplex_13(.clk(clk), .reset(reset),
       .io_real1( fft_5_Y10 ),
       .io_img1( fft_5_Y11 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_13_io_realOut ),
       .io_imgOut( multComplex_13_io_imgOut )
  );
  multComplex multComplex_14(.clk(clk), .reset(reset),
       .io_real1( fft_5_Y12 ),
       .io_img1( fft_5_Y13 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_14_io_realOut ),
       .io_imgOut( multComplex_14_io_imgOut )
  );
  multComplex multComplex_15(.clk(clk), .reset(reset),
       .io_real1( fft_5_Y14 ),
       .io_img1( fft_5_Y15 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_15_io_realOut ),
       .io_imgOut( multComplex_15_io_imgOut )
  );
  multComplex multComplex_16(.clk(clk), .reset(reset),
       .io_real1( fft_6_Y0 ),
       .io_img1( fft_6_Y1 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_16_io_realOut ),
       .io_imgOut( multComplex_16_io_imgOut )
  );
  multComplex multComplex_17(.clk(clk), .reset(reset),
       .io_real1( fft_6_Y2 ),
       .io_img1( fft_6_Y3 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_17_io_realOut ),
       .io_imgOut( multComplex_17_io_imgOut )
  );
  multComplex multComplex_18(.clk(clk), .reset(reset),
       .io_real1( fft_6_Y4 ),
       .io_img1( fft_6_Y5 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_18_io_realOut ),
       .io_imgOut( multComplex_18_io_imgOut )
  );
  multComplex multComplex_19(.clk(clk), .reset(reset),
       .io_real1( fft_6_Y6 ),
       .io_img1( fft_6_Y7 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_19_io_realOut ),
       .io_imgOut( multComplex_19_io_imgOut )
  );
  multComplex multComplex_20(.clk(clk), .reset(reset),
       .io_real1( fft_6_Y8 ),
       .io_img1( fft_6_Y9 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_20_io_realOut ),
       .io_imgOut( multComplex_20_io_imgOut )
  );
  multComplex multComplex_21(.clk(clk), .reset(reset),
       .io_real1( fft_6_Y10 ),
       .io_img1( fft_6_Y11 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_21_io_realOut ),
       .io_imgOut( multComplex_21_io_imgOut )
  );
  multComplex multComplex_22(.clk(clk), .reset(reset),
       .io_real1( fft_6_Y12 ),
       .io_img1( fft_6_Y13 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_22_io_realOut ),
       .io_imgOut( multComplex_22_io_imgOut )
  );
  multComplex multComplex_23(.clk(clk), .reset(reset),
       .io_real1( fft_6_Y14 ),
       .io_img1( fft_6_Y15 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_23_io_realOut ),
       .io_imgOut( multComplex_23_io_imgOut )
  );
  multComplex multComplex_24(.clk(clk), .reset(reset),
       .io_real1( fft_7_Y0 ),
       .io_img1( fft_7_Y1 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_24_io_realOut ),
       .io_imgOut( multComplex_24_io_imgOut )
  );
  multComplex multComplex_25(.clk(clk), .reset(reset),
       .io_real1( fft_7_Y2 ),
       .io_img1( fft_7_Y3 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_25_io_realOut ),
       .io_imgOut( multComplex_25_io_imgOut )
  );
  multComplex multComplex_26(.clk(clk), .reset(reset),
       .io_real1( fft_7_Y4 ),
       .io_img1( fft_7_Y5 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_26_io_realOut ),
       .io_imgOut( multComplex_26_io_imgOut )
  );
  multComplex multComplex_27(.clk(clk), .reset(reset),
       .io_real1( fft_7_Y6 ),
       .io_img1( fft_7_Y7 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_27_io_realOut ),
       .io_imgOut( multComplex_27_io_imgOut )
  );
  multComplex multComplex_28(.clk(clk), .reset(reset),
       .io_real1( fft_7_Y8 ),
       .io_img1( fft_7_Y9 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_28_io_realOut ),
       .io_imgOut( multComplex_28_io_imgOut )
  );
  multComplex multComplex_29(.clk(clk), .reset(reset),
       .io_real1( fft_7_Y10 ),
       .io_img1( fft_7_Y11 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_29_io_realOut ),
       .io_imgOut( multComplex_29_io_imgOut )
  );
  multComplex multComplex_30(.clk(clk), .reset(reset),
       .io_real1( fft_7_Y12 ),
       .io_img1( fft_7_Y13 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_30_io_realOut ),
       .io_imgOut( multComplex_30_io_imgOut )
  );
  multComplex multComplex_31(.clk(clk), .reset(reset),
       .io_real1( fft_7_Y14 ),
       .io_img1( fft_7_Y15 ),
       .io_real2( 16'h1 ),
       .io_img2( 16'h1 ),
       .io_realOut( multComplex_31_io_realOut ),
       .io_imgOut( multComplex_31_io_imgOut )
  );
  ifft8_8 fft_8(.clk(clk), .reset(reset),
       .next( delayArrayNext_2 ),
       .next_out( fft_8_next_out ),
       .X15( multComplex_7_io_imgOut ),
       .X14( multComplex_7_io_realOut ),
       .X13( multComplex_6_io_imgOut ),
       .X12( multComplex_6_io_realOut ),
       .X11( multComplex_5_io_imgOut ),
       .X10( multComplex_5_io_realOut ),
       .X9( multComplex_4_io_imgOut ),
       .X8( multComplex_4_io_realOut ),
       .X7( multComplex_3_io_imgOut ),
       .X6( multComplex_3_io_realOut ),
       .X5( multComplex_2_io_imgOut ),
       .X4( multComplex_2_io_realOut ),
       .X3( multComplex_1_io_imgOut ),
       .X2( multComplex_1_io_realOut ),
       .X1( multComplex_io_imgOut ),
       .X0( multComplex_io_realOut ),
       .Y15( fft_8_Y15 ),
       .Y14( fft_8_Y14 ),
       .Y13( fft_8_Y13 ),
       .Y12( fft_8_Y12 ),
       .Y11( fft_8_Y11 ),
       .Y10( fft_8_Y10 ),
       .Y9( fft_8_Y9 ),
       .Y8( fft_8_Y8 ),
       .Y7( fft_8_Y7 ),
       .Y6( fft_8_Y6 ),
       .Y5( fft_8_Y5 ),
       .Y4( fft_8_Y4 ),
       .Y3( fft_8_Y3 ),
       .Y2( fft_8_Y2 ),
       .Y1( fft_8_Y1 ),
       .Y0( fft_8_Y0 )
  );
  ifft8_8 fft_9(.clk(clk), .reset(reset),
       .next( delayArrayNext_2 ),
       //.next_out(  )
       .X15( multComplex_15_io_imgOut ),
       .X14( multComplex_15_io_realOut ),
       .X13( multComplex_14_io_imgOut ),
       .X12( multComplex_14_io_realOut ),
       .X11( multComplex_13_io_imgOut ),
       .X10( multComplex_13_io_realOut ),
       .X9( multComplex_12_io_imgOut ),
       .X8( multComplex_12_io_realOut ),
       .X7( multComplex_11_io_imgOut ),
       .X6( multComplex_11_io_realOut ),
       .X5( multComplex_10_io_imgOut ),
       .X4( multComplex_10_io_realOut ),
       .X3( multComplex_9_io_imgOut ),
       .X2( multComplex_9_io_realOut ),
       .X1( multComplex_8_io_imgOut ),
       .X0( multComplex_8_io_realOut ),
       .Y15( fft_9_Y15 ),
       .Y14( fft_9_Y14 ),
       .Y13( fft_9_Y13 ),
       .Y12( fft_9_Y12 ),
       .Y11( fft_9_Y11 ),
       .Y10( fft_9_Y10 ),
       .Y9( fft_9_Y9 ),
       .Y8( fft_9_Y8 ),
       .Y7( fft_9_Y7 ),
       .Y6( fft_9_Y6 ),
       .Y5( fft_9_Y5 ),
       .Y4( fft_9_Y4 ),
       .Y3( fft_9_Y3 ),
       .Y2( fft_9_Y2 ),
       .Y1( fft_9_Y1 ),
       .Y0( fft_9_Y0 )
  );
  ifft8_8 fft_10(.clk(clk), .reset(reset),
       .next( delayArrayNext_2 ),
       //.next_out(  )
       .X15( multComplex_23_io_imgOut ),
       .X14( multComplex_23_io_realOut ),
       .X13( multComplex_22_io_imgOut ),
       .X12( multComplex_22_io_realOut ),
       .X11( multComplex_21_io_imgOut ),
       .X10( multComplex_21_io_realOut ),
       .X9( multComplex_20_io_imgOut ),
       .X8( multComplex_20_io_realOut ),
       .X7( multComplex_19_io_imgOut ),
       .X6( multComplex_19_io_realOut ),
       .X5( multComplex_18_io_imgOut ),
       .X4( multComplex_18_io_realOut ),
       .X3( multComplex_17_io_imgOut ),
       .X2( multComplex_17_io_realOut ),
       .X1( multComplex_16_io_imgOut ),
       .X0( multComplex_16_io_realOut ),
       .Y15( fft_10_Y15 ),
       .Y14( fft_10_Y14 ),
       .Y13( fft_10_Y13 ),
       .Y12( fft_10_Y12 ),
       .Y11( fft_10_Y11 ),
       .Y10( fft_10_Y10 ),
       .Y9( fft_10_Y9 ),
       .Y8( fft_10_Y8 ),
       .Y7( fft_10_Y7 ),
       .Y6( fft_10_Y6 ),
       .Y5( fft_10_Y5 ),
       .Y4( fft_10_Y4 ),
       .Y3( fft_10_Y3 ),
       .Y2( fft_10_Y2 ),
       .Y1( fft_10_Y1 ),
       .Y0( fft_10_Y0 )
  );
  ifft8_8 fft_11(.clk(clk), .reset(reset),
       .next( delayArrayNext_2 ),
       //.next_out(  )
       .X15( multComplex_31_io_imgOut ),
       .X14( multComplex_31_io_realOut ),
       .X13( multComplex_30_io_imgOut ),
       .X12( multComplex_30_io_realOut ),
       .X11( multComplex_29_io_imgOut ),
       .X10( multComplex_29_io_realOut ),
       .X9( multComplex_28_io_imgOut ),
       .X8( multComplex_28_io_realOut ),
       .X7( multComplex_27_io_imgOut ),
       .X6( multComplex_27_io_realOut ),
       .X5( multComplex_26_io_imgOut ),
       .X4( multComplex_26_io_realOut ),
       .X3( multComplex_25_io_imgOut ),
       .X2( multComplex_25_io_realOut ),
       .X1( multComplex_24_io_imgOut ),
       .X0( multComplex_24_io_realOut ),
       .Y15( fft_11_Y15 ),
       .Y14( fft_11_Y14 ),
       .Y13( fft_11_Y13 ),
       .Y12( fft_11_Y12 ),
       .Y11( fft_11_Y11 ),
       .Y10( fft_11_Y10 ),
       .Y9( fft_11_Y9 ),
       .Y8( fft_11_Y8 ),
       .Y7( fft_11_Y7 ),
       .Y6( fft_11_Y6 ),
       .Y5( fft_11_Y5 ),
       .Y4( fft_11_Y4 ),
       .Y3( fft_11_Y3 ),
       .Y2( fft_11_Y2 ),
       .Y1( fft_11_Y1 ),
       .Y0( fft_11_Y0 )
  );
  ifft8_8 fft_12(.clk(clk), .reset(reset),
       .next( streamMatrixTransposeTop_1_io_start_next_stage ),
       .next_out( fft_12_next_out ),
       .X15( T95 ),
       .X14( T94 ),
       .X13( T93 ),
       .X12( T92 ),
       .X11( T91 ),
       .X10( T90 ),
       .X9( T89 ),
       .X8( T88 ),
       .X7( T87 ),
       .X6( T86 ),
       .X5( T85 ),
       .X4( T84 ),
       .X3( T83 ),
       .X2( T82 ),
       .X1( T81 ),
       .X0( T80 ),
       //.Y15(  )
       .Y14( fft_12_Y14 ),
       //.Y13(  )
       .Y12( fft_12_Y12 ),
       //.Y11(  )
       .Y10( fft_12_Y10 ),
       //.Y9(  )
       .Y8( fft_12_Y8 ),
       //.Y7(  )
       .Y6( fft_12_Y6 ),
       //.Y5(  )
       .Y4( fft_12_Y4 ),
       //.Y3(  )
       .Y2( fft_12_Y2 ),
       //.Y1(  )
       .Y0( fft_12_Y0 )
  );
  ifft8_8 fft_13(.clk(clk), .reset(reset),
       .next( streamMatrixTransposeTop_1_io_start_next_stage ),
       //.next_out(  )
       .X15( T79 ),
       .X14( T78 ),
       .X13( T77 ),
       .X12( T76 ),
       .X11( T75 ),
       .X10( T74 ),
       .X9( T73 ),
       .X8( T72 ),
       .X7( T71 ),
       .X6( T70 ),
       .X5( T69 ),
       .X4( T68 ),
       .X3( T67 ),
       .X2( T66 ),
       .X1( T65 ),
       .X0( T64 ),
       //.Y15(  )
       .Y14( fft_13_Y14 ),
       //.Y13(  )
       .Y12( fft_13_Y12 ),
       //.Y11(  )
       .Y10( fft_13_Y10 ),
       //.Y9(  )
       .Y8( fft_13_Y8 ),
       //.Y7(  )
       .Y6( fft_13_Y6 ),
       //.Y5(  )
       .Y4( fft_13_Y4 ),
       //.Y3(  )
       .Y2( fft_13_Y2 ),
       //.Y1(  )
       .Y0( fft_13_Y0 )
  );
  ifft8_8 fft_14(.clk(clk), .reset(reset),
       .next( streamMatrixTransposeTop_1_io_start_next_stage ),
       //.next_out(  )
       .X15( T63 ),
       .X14( T62 ),
       .X13( T61 ),
       .X12( T60 ),
       .X11( T59 ),
       .X10( T58 ),
       .X9( T57 ),
       .X8( T56 ),
       .X7( T55 ),
       .X6( T54 ),
       .X5( T53 ),
       .X4( T52 ),
       .X3( T51 ),
       .X2( T50 ),
       .X1( T49 ),
       .X0( T48 ),
       //.Y15(  )
       .Y14( fft_14_Y14 ),
       //.Y13(  )
       .Y12( fft_14_Y12 ),
       //.Y11(  )
       .Y10( fft_14_Y10 ),
       //.Y9(  )
       .Y8( fft_14_Y8 ),
       //.Y7(  )
       .Y6( fft_14_Y6 ),
       //.Y5(  )
       .Y4( fft_14_Y4 ),
       //.Y3(  )
       .Y2( fft_14_Y2 ),
       //.Y1(  )
       .Y0( fft_14_Y0 )
  );
  ifft8_8 fft_15(.clk(clk), .reset(reset),
       .next( streamMatrixTransposeTop_1_io_start_next_stage ),
       //.next_out(  )
       .X15( T47 ),
       .X14( T46 ),
       .X13( T45 ),
       .X12( T44 ),
       .X11( T43 ),
       .X10( T42 ),
       .X9( T41 ),
       .X8( T40 ),
       .X7( T39 ),
       .X6( T38 ),
       .X5( T37 ),
       .X4( T36 ),
       .X3( T35 ),
       .X2( T34 ),
       .X1( T33 ),
       .X0( T32 ),
       //.Y15(  )
       .Y14( fft_15_Y14 ),
       //.Y13(  )
       .Y12( fft_15_Y12 ),
       //.Y11(  )
       .Y10( fft_15_Y10 ),
       //.Y9(  )
       .Y8( fft_15_Y8 ),
       //.Y7(  )
       .Y6( fft_15_Y6 ),
       //.Y5(  )
       .Y4( fft_15_Y4 ),
       //.Y3(  )
       .Y2( fft_15_Y2 ),
       //.Y1(  )
       .Y0( fft_15_Y0 )
  );
  streamMatrixTransposeTop streamMatrixTransposeTop_1(.clk(clk), .reset(reset),
       .io_clk_en( 1'h1 ),
       .io_start( startSecondMatrix ),
       .io_start_next_stage( streamMatrixTransposeTop_1_io_start_next_stage ),
       .io_in_31( T31 ),
       .io_in_30( T30 ),
       .io_in_29( T29 ),
       .io_in_28( T28 ),
       .io_in_27( T27 ),
       .io_in_26( T26 ),
       .io_in_25( T25 ),
       .io_in_24( T24 ),
       .io_in_23( T23 ),
       .io_in_22( T22 ),
       .io_in_21( T21 ),
       .io_in_20( T20 ),
       .io_in_19( T19 ),
       .io_in_18( T18 ),
       .io_in_17( T17 ),
       .io_in_16( T16 ),
       .io_in_15( T15 ),
       .io_in_14( T14 ),
       .io_in_13( T13 ),
       .io_in_12( T12 ),
       .io_in_11( T11 ),
       .io_in_10( T10 ),
       .io_in_9( T9 ),
       .io_in_8( T8 ),
       .io_in_7( T7 ),
       .io_in_6( T6 ),
       .io_in_5( T5 ),
       .io_in_4( T4 ),
       .io_in_3( T3 ),
       .io_in_2( T2 ),
       .io_in_1( T1 ),
       .io_in_0( T0 ),
       .io_out_31( streamMatrixTransposeTop_1_io_out_31 ),
       .io_out_30( streamMatrixTransposeTop_1_io_out_30 ),
       .io_out_29( streamMatrixTransposeTop_1_io_out_29 ),
       .io_out_28( streamMatrixTransposeTop_1_io_out_28 ),
       .io_out_27( streamMatrixTransposeTop_1_io_out_27 ),
       .io_out_26( streamMatrixTransposeTop_1_io_out_26 ),
       .io_out_25( streamMatrixTransposeTop_1_io_out_25 ),
       .io_out_24( streamMatrixTransposeTop_1_io_out_24 ),
       .io_out_23( streamMatrixTransposeTop_1_io_out_23 ),
       .io_out_22( streamMatrixTransposeTop_1_io_out_22 ),
       .io_out_21( streamMatrixTransposeTop_1_io_out_21 ),
       .io_out_20( streamMatrixTransposeTop_1_io_out_20 ),
       .io_out_19( streamMatrixTransposeTop_1_io_out_19 ),
       .io_out_18( streamMatrixTransposeTop_1_io_out_18 ),
       .io_out_17( streamMatrixTransposeTop_1_io_out_17 ),
       .io_out_16( streamMatrixTransposeTop_1_io_out_16 ),
       .io_out_15( streamMatrixTransposeTop_1_io_out_15 ),
       .io_out_14( streamMatrixTransposeTop_1_io_out_14 ),
       .io_out_13( streamMatrixTransposeTop_1_io_out_13 ),
       .io_out_12( streamMatrixTransposeTop_1_io_out_12 ),
       .io_out_11( streamMatrixTransposeTop_1_io_out_11 ),
       .io_out_10( streamMatrixTransposeTop_1_io_out_10 ),
       .io_out_9( streamMatrixTransposeTop_1_io_out_9 ),
       .io_out_8( streamMatrixTransposeTop_1_io_out_8 ),
       .io_out_7( streamMatrixTransposeTop_1_io_out_7 ),
       .io_out_6( streamMatrixTransposeTop_1_io_out_6 ),
       .io_out_5( streamMatrixTransposeTop_1_io_out_5 ),
       .io_out_4( streamMatrixTransposeTop_1_io_out_4 ),
       .io_out_3( streamMatrixTransposeTop_1_io_out_3 ),
       .io_out_2( streamMatrixTransposeTop_1_io_out_2 ),
       .io_out_1( streamMatrixTransposeTop_1_io_out_1 ),
       .io_out_0( streamMatrixTransposeTop_1_io_out_0 )
  );

  always @(posedge clk) begin
    startSecondMatrix <= fft_8_next_out;
    delaySecond_24 <= streamMatrixTransposeTop_1_io_out_24;
    delaySecond_25 <= streamMatrixTransposeTop_1_io_out_25;
    delaySecond_26 <= streamMatrixTransposeTop_1_io_out_26;
    delaySecond_27 <= streamMatrixTransposeTop_1_io_out_27;
    delaySecond_28 <= streamMatrixTransposeTop_1_io_out_28;
    delaySecond_29 <= streamMatrixTransposeTop_1_io_out_29;
    delaySecond_30 <= streamMatrixTransposeTop_1_io_out_30;
    delaySecond_31 <= streamMatrixTransposeTop_1_io_out_31;
    delaySecond_16 <= streamMatrixTransposeTop_1_io_out_16;
    delaySecond_17 <= streamMatrixTransposeTop_1_io_out_17;
    delaySecond_18 <= streamMatrixTransposeTop_1_io_out_18;
    delaySecond_19 <= streamMatrixTransposeTop_1_io_out_19;
    delaySecond_20 <= streamMatrixTransposeTop_1_io_out_20;
    delaySecond_21 <= streamMatrixTransposeTop_1_io_out_21;
    delaySecond_22 <= streamMatrixTransposeTop_1_io_out_22;
    delaySecond_23 <= streamMatrixTransposeTop_1_io_out_23;
    delaySecond_8 <= streamMatrixTransposeTop_1_io_out_8;
    delaySecond_9 <= streamMatrixTransposeTop_1_io_out_9;
    delaySecond_10 <= streamMatrixTransposeTop_1_io_out_10;
    delaySecond_11 <= streamMatrixTransposeTop_1_io_out_11;
    delaySecond_12 <= streamMatrixTransposeTop_1_io_out_12;
    delaySecond_13 <= streamMatrixTransposeTop_1_io_out_13;
    delaySecond_14 <= streamMatrixTransposeTop_1_io_out_14;
    delaySecond_15 <= streamMatrixTransposeTop_1_io_out_15;
    delaySecond_0 <= streamMatrixTransposeTop_1_io_out_0;
    delaySecond_1 <= streamMatrixTransposeTop_1_io_out_1;
    delaySecond_2 <= streamMatrixTransposeTop_1_io_out_2;
    delaySecond_3 <= streamMatrixTransposeTop_1_io_out_3;
    delaySecond_4 <= streamMatrixTransposeTop_1_io_out_4;
    delaySecond_5 <= streamMatrixTransposeTop_1_io_out_5;
    delaySecond_6 <= streamMatrixTransposeTop_1_io_out_6;
    delaySecond_7 <= streamMatrixTransposeTop_1_io_out_7;
    delayArrayNext_2 <= delayArrayNext_1;
    delayArrayNext_1 <= delayArrayNext_0;
    delayArrayNext_0 <= fft_4_next_out;
    delayFirst_24 <= streamMatrixTransposeTop_io_out_24;
    delayFirst_25 <= streamMatrixTransposeTop_io_out_25;
    delayFirst_26 <= streamMatrixTransposeTop_io_out_26;
    delayFirst_27 <= streamMatrixTransposeTop_io_out_27;
    delayFirst_28 <= streamMatrixTransposeTop_io_out_28;
    delayFirst_29 <= streamMatrixTransposeTop_io_out_29;
    delayFirst_30 <= streamMatrixTransposeTop_io_out_30;
    delayFirst_31 <= streamMatrixTransposeTop_io_out_31;
    delayFirst_16 <= streamMatrixTransposeTop_io_out_16;
    delayFirst_17 <= streamMatrixTransposeTop_io_out_17;
    delayFirst_18 <= streamMatrixTransposeTop_io_out_18;
    delayFirst_19 <= streamMatrixTransposeTop_io_out_19;
    delayFirst_20 <= streamMatrixTransposeTop_io_out_20;
    delayFirst_21 <= streamMatrixTransposeTop_io_out_21;
    delayFirst_22 <= streamMatrixTransposeTop_io_out_22;
    delayFirst_23 <= streamMatrixTransposeTop_io_out_23;
    delayFirst_8 <= streamMatrixTransposeTop_io_out_8;
    delayFirst_9 <= streamMatrixTransposeTop_io_out_9;
    delayFirst_10 <= streamMatrixTransposeTop_io_out_10;
    delayFirst_11 <= streamMatrixTransposeTop_io_out_11;
    delayFirst_12 <= streamMatrixTransposeTop_io_out_12;
    delayFirst_13 <= streamMatrixTransposeTop_io_out_13;
    delayFirst_14 <= streamMatrixTransposeTop_io_out_14;
    delayFirst_15 <= streamMatrixTransposeTop_io_out_15;
    delayFirst_0 <= streamMatrixTransposeTop_io_out_0;
    delayFirst_1 <= streamMatrixTransposeTop_io_out_1;
    delayFirst_2 <= streamMatrixTransposeTop_io_out_2;
    delayFirst_3 <= streamMatrixTransposeTop_io_out_3;
    delayFirst_4 <= streamMatrixTransposeTop_io_out_4;
    delayFirst_5 <= streamMatrixTransposeTop_io_out_5;
    delayFirst_6 <= streamMatrixTransposeTop_io_out_6;
    delayFirst_7 <= streamMatrixTransposeTop_io_out_7;
    startFirstMatrix <= fft_next_out;
    delayInput_24 <= io_in_24;
    delayInput_25 <= io_in_25;
    delayInput_26 <= io_in_26;
    delayInput_27 <= io_in_27;
    delayInput_28 <= io_in_28;
    delayInput_29 <= io_in_29;
    delayInput_30 <= io_in_30;
    delayInput_31 <= io_in_31;
    delayInput_16 <= io_in_16;
    delayInput_17 <= io_in_17;
    delayInput_18 <= io_in_18;
    delayInput_19 <= io_in_19;
    delayInput_20 <= io_in_20;
    delayInput_21 <= io_in_21;
    delayInput_22 <= io_in_22;
    delayInput_23 <= io_in_23;
    delayInput_8 <= io_in_8;
    delayInput_9 <= io_in_9;
    delayInput_10 <= io_in_10;
    delayInput_11 <= io_in_11;
    delayInput_12 <= io_in_12;
    delayInput_13 <= io_in_13;
    delayInput_14 <= io_in_14;
    delayInput_15 <= io_in_15;
    delayInput_0 <= io_in_0;
    delayInput_1 <= io_in_1;
    delayInput_2 <= io_in_2;
    delayInput_3 <= io_in_3;
    delayInput_4 <= io_in_4;
    delayInput_5 <= io_in_5;
    delayInput_6 <= io_in_6;
    delayInput_7 <= io_in_7;
    delayStartNextStage <= fft_12_next_out;
  end
endmodule

module afu_user(input clk, input reset,
    input [511:0] input_fifo_din,
    input  input_fifo_we,
    output input_fifo_full,
    output input_fifo_almost_full,
    output[5:0] input_fifo_count,
    output[511:0] output_fifo_dout,
    input  output_fifo_re,
    output output_fifo_empty,
    output output_fifo_almost_empty,
    input [31:0] ctx_length
);

  wire T0;
  wire T1;
  wire T2;
  reg [31:0] ctx_output_count;
  wire[31:0] T90;
  wire[31:0] T3;
  wire[31:0] T4;
  wire[511:0] T5;
  wire[511:0] T6;
  wire[511:0] T7;
  wire[255:0] T8;
  wire[127:0] T9;
  wire[63:0] T10;
  wire[31:0] T11;
  wire[31:0] T12;
  wire[63:0] T13;
  wire[31:0] T14;
  wire[31:0] T15;
  wire[127:0] T16;
  wire[63:0] T17;
  wire[31:0] T18;
  wire[31:0] T19;
  wire[63:0] T20;
  wire[31:0] T21;
  wire[31:0] T22;
  wire[255:0] T23;
  wire[127:0] T24;
  wire[63:0] T25;
  wire[31:0] T26;
  wire[31:0] T27;
  wire[63:0] T28;
  wire[31:0] T29;
  wire[31:0] T30;
  wire[127:0] T31;
  wire[63:0] T32;
  wire[31:0] T33;
  wire[31:0] T34;
  wire[63:0] T35;
  wire[31:0] T36;
  wire[31:0] T37;
  wire[511:0] T38;
  reg [31:0] total_time_count;
  wire[31:0] T91;
  wire[31:0] T39;
  wire[31:0] T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  reg  state;
  wire T92;
  wire T45;
  wire T46;
  wire T47;
  wire[31:0] T48;
  wire[15:0] T49;
  wire[15:0] T50;
  wire[15:0] T51;
  wire[15:0] T52;
  wire[15:0] T53;
  wire[15:0] T54;
  wire[15:0] T55;
  wire[15:0] T56;
  wire[15:0] T57;
  wire[15:0] T58;
  wire[15:0] T59;
  wire[15:0] T60;
  wire[15:0] T61;
  wire[15:0] T62;
  wire[15:0] T63;
  wire[15:0] T64;
  wire[15:0] T65;
  wire[15:0] T66;
  wire[15:0] T67;
  wire[15:0] T68;
  wire[15:0] T69;
  wire[15:0] T70;
  wire[15:0] T71;
  wire[15:0] T72;
  wire[15:0] T73;
  wire[15:0] T74;
  wire[15:0] T75;
  wire[15:0] T76;
  wire[15:0] T77;
  wire[15:0] T78;
  wire[15:0] T79;
  wire[15:0] T80;
  reg  start_reg;
  wire T93;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  reg [31:0] ctx_input_count;
  wire[31:0] T94;
  wire[31:0] T86;
  wire[31:0] T87;
  wire T88;
  wire T89;
  wire[5:0] T95;
  wire[511:0] syn_read_fifo_dout;
  wire syn_read_fifo_empty;
  wire syn_read_fifo_full;
  wire syn_read_fifo_count;
  wire syn_read_fifo_almostfull;
  wire[511:0] syn_read_fifo_1_dout;
  wire syn_read_fifo_1_empty;
  wire syn_read_fifo_1_almostempty;
  wire two_d_convolution_io_start_next_stage;
  wire[15:0] two_d_convolution_io_out_31;
  wire[15:0] two_d_convolution_io_out_30;
  wire[15:0] two_d_convolution_io_out_29;
  wire[15:0] two_d_convolution_io_out_28;
  wire[15:0] two_d_convolution_io_out_27;
  wire[15:0] two_d_convolution_io_out_26;
  wire[15:0] two_d_convolution_io_out_25;
  wire[15:0] two_d_convolution_io_out_24;
  wire[15:0] two_d_convolution_io_out_23;
  wire[15:0] two_d_convolution_io_out_22;
  wire[15:0] two_d_convolution_io_out_21;
  wire[15:0] two_d_convolution_io_out_20;
  wire[15:0] two_d_convolution_io_out_19;
  wire[15:0] two_d_convolution_io_out_18;
  wire[15:0] two_d_convolution_io_out_17;
  wire[15:0] two_d_convolution_io_out_16;
  wire[15:0] two_d_convolution_io_out_15;
  wire[15:0] two_d_convolution_io_out_14;
  wire[15:0] two_d_convolution_io_out_13;
  wire[15:0] two_d_convolution_io_out_12;
  wire[15:0] two_d_convolution_io_out_11;
  wire[15:0] two_d_convolution_io_out_10;
  wire[15:0] two_d_convolution_io_out_9;
  wire[15:0] two_d_convolution_io_out_8;
  wire[15:0] two_d_convolution_io_out_7;
  wire[15:0] two_d_convolution_io_out_6;
  wire[15:0] two_d_convolution_io_out_5;
  wire[15:0] two_d_convolution_io_out_4;
  wire[15:0] two_d_convolution_io_out_3;
  wire[15:0] two_d_convolution_io_out_2;
  wire[15:0] two_d_convolution_io_out_1;
  wire[15:0] two_d_convolution_io_out_0;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    ctx_output_count = {1{$random}};
    total_time_count = {1{$random}};
    state = {1{$random}};
    start_reg = {1{$random}};
    ctx_input_count = {1{$random}};
  end
// synthesis translate_on
`endif

  assign T0 = T2 ? 1'h0 : T1;
  assign T1 = two_d_convolution_io_start_next_stage & T84;
  assign T2 = ctx_length == ctx_output_count;
  assign T90 = reset ? 32'h0 : T3;
  assign T3 = T0 ? T4 : ctx_output_count;
  assign T4 = ctx_output_count + 32'h1;
  assign T5 = T47 ? T38 : T6;
  assign T6 = T7;
  assign T7 = {T23, T8};
  assign T8 = {T16, T9};
  assign T9 = {T13, T10};
  assign T10 = {T12, T11};
  assign T11 = {two_d_convolution_io_out_1, two_d_convolution_io_out_0};
  assign T12 = {two_d_convolution_io_out_3, two_d_convolution_io_out_2};
  assign T13 = {T15, T14};
  assign T14 = {two_d_convolution_io_out_5, two_d_convolution_io_out_4};
  assign T15 = {two_d_convolution_io_out_7, two_d_convolution_io_out_6};
  assign T16 = {T20, T17};
  assign T17 = {T19, T18};
  assign T18 = {two_d_convolution_io_out_9, two_d_convolution_io_out_8};
  assign T19 = {two_d_convolution_io_out_11, two_d_convolution_io_out_10};
  assign T20 = {T22, T21};
  assign T21 = {two_d_convolution_io_out_13, two_d_convolution_io_out_12};
  assign T22 = {two_d_convolution_io_out_15, two_d_convolution_io_out_14};
  assign T23 = {T31, T24};
  assign T24 = {T28, T25};
  assign T25 = {T27, T26};
  assign T26 = {two_d_convolution_io_out_17, two_d_convolution_io_out_16};
  assign T27 = {two_d_convolution_io_out_19, two_d_convolution_io_out_18};
  assign T28 = {T30, T29};
  assign T29 = {two_d_convolution_io_out_21, two_d_convolution_io_out_20};
  assign T30 = {two_d_convolution_io_out_23, two_d_convolution_io_out_22};
  assign T31 = {T35, T32};
  assign T32 = {T34, T33};
  assign T33 = {two_d_convolution_io_out_25, two_d_convolution_io_out_24};
  assign T34 = {two_d_convolution_io_out_27, two_d_convolution_io_out_26};
  assign T35 = {T37, T36};
  assign T36 = {two_d_convolution_io_out_29, two_d_convolution_io_out_28};
  assign T37 = {two_d_convolution_io_out_31, two_d_convolution_io_out_30};
  assign T38 = {480'h0, total_time_count};
  assign T91 = reset ? 32'h0 : T39;
  assign T39 = T41 ? T40 : total_time_count;
  assign T40 = total_time_count + 32'h1;
  assign T41 = T43 & T42;
  assign T42 = ctx_output_count != ctx_length;
  assign T43 = T44 ^ 1'h1;
  assign T44 = state == 1'h0;
  assign T92 = reset ? 1'h0 : T45;
  assign T45 = T46 ? 1'h1 : state;
  assign T46 = T44 & T0;
  assign T47 = T48 == ctx_output_count;
  assign T48 = ctx_length - 32'h1;
  assign T49 = syn_read_fifo_dout[15:0];
  assign T50 = syn_read_fifo_dout[31:16];
  assign T51 = syn_read_fifo_dout[47:32];
  assign T52 = syn_read_fifo_dout[63:48];
  assign T53 = syn_read_fifo_dout[79:64];
  assign T54 = syn_read_fifo_dout[95:80];
  assign T55 = syn_read_fifo_dout[111:96];
  assign T56 = syn_read_fifo_dout[127:112];
  assign T57 = syn_read_fifo_dout[143:128];
  assign T58 = syn_read_fifo_dout[159:144];
  assign T59 = syn_read_fifo_dout[175:160];
  assign T60 = syn_read_fifo_dout[191:176];
  assign T61 = syn_read_fifo_dout[207:192];
  assign T62 = syn_read_fifo_dout[223:208];
  assign T63 = syn_read_fifo_dout[239:224];
  assign T64 = syn_read_fifo_dout[255:240];
  assign T65 = syn_read_fifo_dout[271:256];
  assign T66 = syn_read_fifo_dout[287:272];
  assign T67 = syn_read_fifo_dout[303:288];
  assign T68 = syn_read_fifo_dout[319:304];
  assign T69 = syn_read_fifo_dout[335:320];
  assign T70 = syn_read_fifo_dout[351:336];
  assign T71 = syn_read_fifo_dout[367:352];
  assign T72 = syn_read_fifo_dout[383:368];
  assign T73 = syn_read_fifo_dout[399:384];
  assign T74 = syn_read_fifo_dout[415:400];
  assign T75 = syn_read_fifo_dout[431:416];
  assign T76 = syn_read_fifo_dout[447:432];
  assign T77 = syn_read_fifo_dout[463:448];
  assign T78 = syn_read_fifo_dout[479:464];
  assign T79 = syn_read_fifo_dout[495:480];
  assign T80 = syn_read_fifo_dout[511:496];
  assign T93 = reset ? 1'h0 : T81;
  assign T81 = T83 ? 1'h0 : T82;
  assign T82 = T88 ? 1'h1 : start_reg;
  assign T83 = T88 ^ 1'h1;
  assign T84 = T85 ? 1'h1 : start_reg;
  assign T85 = ctx_length == ctx_input_count;
  assign T94 = reset ? 32'h0 : T86;
  assign T86 = T88 ? T87 : ctx_input_count;
  assign T87 = ctx_input_count + 32'h1;
  assign T88 = reset ? 1'h0 : T89;
  assign T89 = ~ syn_read_fifo_empty;
  assign output_fifo_almost_empty = syn_read_fifo_1_almostempty;
  assign output_fifo_empty = syn_read_fifo_1_empty;
  assign output_fifo_dout = syn_read_fifo_1_dout;
  assign input_fifo_count = T95;
  assign T95 = {5'h0, syn_read_fifo_count};
  assign input_fifo_almost_full = syn_read_fifo_almostfull;
  assign input_fifo_full = syn_read_fifo_full;
  syn_read_fifo #(.FIFO_WIDTH(512),.FIFO_DEPTH_BITS(6),.FIFO_ALMOSTFULL_THRESHOLD(60),.FIFO_ALMOSTEMPTY_THRESHOLD(2))
  syn_read_fifo(.clk(clk), .reset(reset),
       .din( input_fifo_din ),
       .we( input_fifo_we ),
       .re( T88 ),
       .dout( syn_read_fifo_dout ),
       .empty( syn_read_fifo_empty ),
       //.almostempty(  )
       .full( syn_read_fifo_full ),
       .count( syn_read_fifo_count ),
       .almostfull( syn_read_fifo_almostfull )
  );
  two_d_convolution two_d_convolution(.clk(clk), .reset(reset),
       .io_clk_en( T84 ),
       .io_start( start_reg ),
       .io_start_next_stage( two_d_convolution_io_start_next_stage ),
       .io_in_31( T80 ),
       .io_in_30( T79 ),
       .io_in_29( T78 ),
       .io_in_28( T77 ),
       .io_in_27( T76 ),
       .io_in_26( T75 ),
       .io_in_25( T74 ),
       .io_in_24( T73 ),
       .io_in_23( T72 ),
       .io_in_22( T71 ),
       .io_in_21( T70 ),
       .io_in_20( T69 ),
       .io_in_19( T68 ),
       .io_in_18( T67 ),
       .io_in_17( T66 ),
       .io_in_16( T65 ),
       .io_in_15( T64 ),
       .io_in_14( T63 ),
       .io_in_13( T62 ),
       .io_in_12( T61 ),
       .io_in_11( T60 ),
       .io_in_10( T59 ),
       .io_in_9( T58 ),
       .io_in_8( T57 ),
       .io_in_7( T56 ),
       .io_in_6( T55 ),
       .io_in_5( T54 ),
       .io_in_4( T53 ),
       .io_in_3( T52 ),
       .io_in_2( T51 ),
       .io_in_1( T50 ),
       .io_in_0( T49 ),
       .io_out_31( two_d_convolution_io_out_31 ),
       .io_out_30( two_d_convolution_io_out_30 ),
       .io_out_29( two_d_convolution_io_out_29 ),
       .io_out_28( two_d_convolution_io_out_28 ),
       .io_out_27( two_d_convolution_io_out_27 ),
       .io_out_26( two_d_convolution_io_out_26 ),
       .io_out_25( two_d_convolution_io_out_25 ),
       .io_out_24( two_d_convolution_io_out_24 ),
       .io_out_23( two_d_convolution_io_out_23 ),
       .io_out_22( two_d_convolution_io_out_22 ),
       .io_out_21( two_d_convolution_io_out_21 ),
       .io_out_20( two_d_convolution_io_out_20 ),
       .io_out_19( two_d_convolution_io_out_19 ),
       .io_out_18( two_d_convolution_io_out_18 ),
       .io_out_17( two_d_convolution_io_out_17 ),
       .io_out_16( two_d_convolution_io_out_16 ),
       .io_out_15( two_d_convolution_io_out_15 ),
       .io_out_14( two_d_convolution_io_out_14 ),
       .io_out_13( two_d_convolution_io_out_13 ),
       .io_out_12( two_d_convolution_io_out_12 ),
       .io_out_11( two_d_convolution_io_out_11 ),
       .io_out_10( two_d_convolution_io_out_10 ),
       .io_out_9( two_d_convolution_io_out_9 ),
       .io_out_8( two_d_convolution_io_out_8 ),
       .io_out_7( two_d_convolution_io_out_7 ),
       .io_out_6( two_d_convolution_io_out_6 ),
       .io_out_5( two_d_convolution_io_out_5 ),
       .io_out_4( two_d_convolution_io_out_4 ),
       .io_out_3( two_d_convolution_io_out_3 ),
       .io_out_2( two_d_convolution_io_out_2 ),
       .io_out_1( two_d_convolution_io_out_1 ),
       .io_out_0( two_d_convolution_io_out_0 )
  );
  syn_read_fifo #(.FIFO_WIDTH(512),.FIFO_DEPTH_BITS(6),.FIFO_ALMOSTFULL_THRESHOLD(60),.FIFO_ALMOSTEMPTY_THRESHOLD(2))
  syn_read_fifo_1(.clk(clk), .reset(reset),
       .din( T5 ),
       .we( T0 ),
       .re( output_fifo_re ),
       .dout( syn_read_fifo_1_dout ),
       .empty( syn_read_fifo_1_empty ),
       .almostempty( syn_read_fifo_1_almostempty )
       //.full(  )
       //.count(  )
       //.almostfull(  )
  );

  always @(posedge clk) begin
    if(reset) begin
      ctx_output_count <= 32'h0;
    end else if(T0) begin
      ctx_output_count <= T4;
    end
    if(reset) begin
      total_time_count <= 32'h0;
    end else if(T41) begin
      total_time_count <= T40;
    end
    if(reset) begin
      state <= 1'h0;
    end else if(T46) begin
      state <= 1'h1;
    end
    if(reset) begin
      start_reg <= 1'h0;
    end else if(T83) begin
      start_reg <= 1'h0;
    end else if(T88) begin
      start_reg <= 1'h1;
    end
    if(reset) begin
      ctx_input_count <= 32'h0;
    end else if(T88) begin
      ctx_input_count <= T87;
    end
  end
endmodule

